-- Banco de pruebas de Tabla de consulta de Datos
-- 
-- Diseño Lógico
-- Gustavo David Mendoza Pinto

LIBRARY IEEE; 
USE IEEE.std_logic_1164.all; 
Entity TB_binary_SevenSegments is 
	
END TB_binary_SevenSegments; 
Architecture Simulation of TB_binary_SevenSegments is 
	Component binary_SevenSegments
		 port(
			 X : in  std_logic_vector(7 downto 0);
			 Y : out std_logic_vector(27 downto 0));
	end Component; 
	 signal X : std_logic_vector(7 downto 0);
	 signal Y : std_logic_vector(27 downto 0)
;BEGIN 
		 SIMBLK00: binary_SevenSegments PORT MAP(X,Y);
	 process 
	 begin 
			 X <="00000000";
			 wait for 20 ns;
			 X <="00000001";
			 wait for 20 ns;
			 X <="00000010";
			 wait for 20 ns;
			 X <="00000011";
			 wait for 20 ns;
			 X <="00000100";
			 wait for 20 ns;
			 X <="00000101";
			 wait for 20 ns;
			 X <="00000110";
			 wait for 20 ns;
			 X <="00000111";
			 wait for 20 ns;
			 X <="00001000";
			 wait for 20 ns;
			 X <="00001001";
			 wait for 20 ns;
			 X <="00001010";
			 wait for 20 ns;
			 X <="00001011";
			 wait for 20 ns;
			 X <="00001100";
			 wait for 20 ns;
			 X <="00001101";
			 wait for 20 ns;
			 X <="00001110";
			 wait for 20 ns;
			 X <="00001111";
			 wait for 20 ns;
			 X <="00010000";
			 wait for 20 ns;
			 X <="00010001";
			 wait for 20 ns;
			 X <="00010010";
			 wait for 20 ns;
			 X <="00010011";
			 wait for 20 ns;
			 X <="00010100";
			 wait for 20 ns;
			 X <="00010101";
			 wait for 20 ns;
			 X <="00010110";
			 wait for 20 ns;
			 X <="00010111";
			 wait for 20 ns;
			 X <="00011000";
			 wait for 20 ns;
			 X <="00011001";
			 wait for 20 ns;
			 X <="00011010";
			 wait for 20 ns;
			 X <="00011011";
			 wait for 20 ns;
			 X <="00011100";
			 wait for 20 ns;
			 X <="00011101";
			 wait for 20 ns;
			 X <="00011110";
			 wait for 20 ns;
			 X <="00011111";
			 wait for 20 ns;
			 X <="00100000";
			 wait for 20 ns;
			 X <="00100001";
			 wait for 20 ns;
			 X <="00100010";
			 wait for 20 ns;
			 X <="00100011";
			 wait for 20 ns;
			 X <="00100100";
			 wait for 20 ns;
			 X <="00100101";
			 wait for 20 ns;
			 X <="00100110";
			 wait for 20 ns;
			 X <="00100111";
			 wait for 20 ns;
			 X <="00101000";
			 wait for 20 ns;
			 X <="00101001";
			 wait for 20 ns;
			 X <="00101010";
			 wait for 20 ns;
			 X <="00101011";
			 wait for 20 ns;
			 X <="00101100";
			 wait for 20 ns;
			 X <="00101101";
			 wait for 20 ns;
			 X <="00101110";
			 wait for 20 ns;
			 X <="00101111";
			 wait for 20 ns;
			 X <="00110000";
			 wait for 20 ns;
			 X <="00110001";
			 wait for 20 ns;
			 X <="00110010";
			 wait for 20 ns;
			 X <="00110011";
			 wait for 20 ns;
			 X <="00110100";
			 wait for 20 ns;
			 X <="00110101";
			 wait for 20 ns;
			 X <="00110110";
			 wait for 20 ns;
			 X <="00110111";
			 wait for 20 ns;
			 X <="00111000";
			 wait for 20 ns;
			 X <="00111001";
			 wait for 20 ns;
			 X <="00111010";
			 wait for 20 ns;
			 X <="00111011";
			 wait for 20 ns;
			 X <="00111100";
			 wait for 20 ns;
			 X <="00111101";
			 wait for 20 ns;
			 X <="00111110";
			 wait for 20 ns;
			 X <="00111111";
			 wait for 20 ns;
			 X <="01000000";
			 wait for 20 ns;
			 X <="01000001";
			 wait for 20 ns;
			 X <="01000010";
			 wait for 20 ns;
			 X <="01000011";
			 wait for 20 ns;
			 X <="01000100";
			 wait for 20 ns;
			 X <="01000101";
			 wait for 20 ns;
			 X <="01000110";
			 wait for 20 ns;
			 X <="01000111";
			 wait for 20 ns;
			 X <="01001000";
			 wait for 20 ns;
			 X <="01001001";
			 wait for 20 ns;
			 X <="01001010";
			 wait for 20 ns;
			 X <="01001011";
			 wait for 20 ns;
			 X <="01001100";
			 wait for 20 ns;
			 X <="01001101";
			 wait for 20 ns;
			 X <="01001110";
			 wait for 20 ns;
			 X <="01001111";
			 wait for 20 ns;
			 X <="01010000";
			 wait for 20 ns;
			 X <="01010001";
			 wait for 20 ns;
			 X <="01010010";
			 wait for 20 ns;
			 X <="01010011";
			 wait for 20 ns;
			 X <="01010100";
			 wait for 20 ns;
			 X <="01010101";
			 wait for 20 ns;
			 X <="01010110";
			 wait for 20 ns;
			 X <="01010111";
			 wait for 20 ns;
			 X <="01011000";
			 wait for 20 ns;
			 X <="01011001";
			 wait for 20 ns;
			 X <="01011010";
			 wait for 20 ns;
			 X <="01011011";
			 wait for 20 ns;
			 X <="01011100";
			 wait for 20 ns;
			 X <="01011101";
			 wait for 20 ns;
			 X <="01011110";
			 wait for 20 ns;
			 X <="01011111";
			 wait for 20 ns;
			 X <="01100000";
			 wait for 20 ns;
			 X <="01100001";
			 wait for 20 ns;
			 X <="01100010";
			 wait for 20 ns;
			 X <="01100011";
			 wait for 20 ns;
			 X <="01100100";
			 wait for 20 ns;
			 X <="01100101";
			 wait for 20 ns;
			 X <="01100110";
			 wait for 20 ns;
			 X <="01100111";
			 wait for 20 ns;
			 X <="01101000";
			 wait for 20 ns;
			 X <="01101001";
			 wait for 20 ns;
			 X <="01101010";
			 wait for 20 ns;
			 X <="01101011";
			 wait for 20 ns;
			 X <="01101100";
			 wait for 20 ns;
			 X <="01101101";
			 wait for 20 ns;
			 X <="01101110";
			 wait for 20 ns;
			 X <="01101111";
			 wait for 20 ns;
			 X <="01110000";
			 wait for 20 ns;
			 X <="01110001";
			 wait for 20 ns;
			 X <="01110010";
			 wait for 20 ns;
			 X <="01110011";
			 wait for 20 ns;
			 X <="01110100";
			 wait for 20 ns;
			 X <="01110101";
			 wait for 20 ns;
			 X <="01110110";
			 wait for 20 ns;
			 X <="01110111";
			 wait for 20 ns;
			 X <="01111000";
			 wait for 20 ns;
			 X <="01111001";
			 wait for 20 ns;
			 X <="01111010";
			 wait for 20 ns;
			 X <="01111011";
			 wait for 20 ns;
			 X <="01111100";
			 wait for 20 ns;
			 X <="01111101";
			 wait for 20 ns;
			 X <="01111110";
			 wait for 20 ns;
			 X <="01111111";
			 wait for 20 ns;
			 X <="10000000";
			 wait for 20 ns;
			 X <="10000001";
			 wait for 20 ns;
			 X <="10000010";
			 wait for 20 ns;
			 X <="10000011";
			 wait for 20 ns;
			 X <="10000100";
			 wait for 20 ns;
			 X <="10000101";
			 wait for 20 ns;
			 X <="10000110";
			 wait for 20 ns;
			 X <="10000111";
			 wait for 20 ns;
			 X <="10001000";
			 wait for 20 ns;
			 X <="10001001";
			 wait for 20 ns;
			 X <="10001010";
			 wait for 20 ns;
			 X <="10001011";
			 wait for 20 ns;
			 X <="10001100";
			 wait for 20 ns;
			 X <="10001101";
			 wait for 20 ns;
			 X <="10001110";
			 wait for 20 ns;
			 X <="10001111";
			 wait for 20 ns;
			 X <="10010000";
			 wait for 20 ns;
			 X <="10010001";
			 wait for 20 ns;
			 X <="10010010";
			 wait for 20 ns;
			 X <="10010011";
			 wait for 20 ns;
			 X <="10010100";
			 wait for 20 ns;
			 X <="10010101";
			 wait for 20 ns;
			 X <="10010110";
			 wait for 20 ns;
			 X <="10010111";
			 wait for 20 ns;
			 X <="10011000";
			 wait for 20 ns;
			 X <="10011001";
			 wait for 20 ns;
			 X <="10011010";
			 wait for 20 ns;
			 X <="10011011";
			 wait for 20 ns;
			 X <="10011100";
			 wait for 20 ns;
			 X <="10011101";
			 wait for 20 ns;
			 X <="10011110";
			 wait for 20 ns;
			 X <="10011111";
			 wait for 20 ns;
			 X <="10100000";
			 wait for 20 ns;
			 X <="10100001";
			 wait for 20 ns;
			 X <="10100010";
			 wait for 20 ns;
			 X <="10100011";
			 wait for 20 ns;
			 X <="10100100";
			 wait for 20 ns;
			 X <="10100101";
			 wait for 20 ns;
			 X <="10100110";
			 wait for 20 ns;
			 X <="10100111";
			 wait for 20 ns;
			 X <="10101000";
			 wait for 20 ns;
			 X <="10101001";
			 wait for 20 ns;
			 X <="10101010";
			 wait for 20 ns;
			 X <="10101011";
			 wait for 20 ns;
			 X <="10101100";
			 wait for 20 ns;
			 X <="10101101";
			 wait for 20 ns;
			 X <="10101110";
			 wait for 20 ns;
			 X <="10101111";
			 wait for 20 ns;
			 X <="10110000";
			 wait for 20 ns;
			 X <="10110001";
			 wait for 20 ns;
			 X <="10110010";
			 wait for 20 ns;
			 X <="10110011";
			 wait for 20 ns;
			 X <="10110100";
			 wait for 20 ns;
			 X <="10110101";
			 wait for 20 ns;
			 X <="10110110";
			 wait for 20 ns;
			 X <="10110111";
			 wait for 20 ns;
			 X <="10111000";
			 wait for 20 ns;
			 X <="10111001";
			 wait for 20 ns;
			 X <="10111010";
			 wait for 20 ns;
			 X <="10111011";
			 wait for 20 ns;
			 X <="10111100";
			 wait for 20 ns;
			 X <="10111101";
			 wait for 20 ns;
			 X <="10111110";
			 wait for 20 ns;
			 X <="10111111";
			 wait for 20 ns;
			 X <="11000000";
			 wait for 20 ns;
			 X <="11000001";
			 wait for 20 ns;
			 X <="11000010";
			 wait for 20 ns;
			 X <="11000011";
			 wait for 20 ns;
			 X <="11000100";
			 wait for 20 ns;
			 X <="11000101";
			 wait for 20 ns;
			 X <="11000110";
			 wait for 20 ns;
			 X <="11000111";
			 wait for 20 ns;
			 X <="11001000";
			 wait for 20 ns;
			 X <="11001001";
			 wait for 20 ns;
			 X <="11001010";
			 wait for 20 ns;
			 X <="11001011";
			 wait for 20 ns;
			 X <="11001100";
			 wait for 20 ns;
			 X <="11001101";
			 wait for 20 ns;
			 X <="11001110";
			 wait for 20 ns;
			 X <="11001111";
			 wait for 20 ns;
			 X <="11010000";
			 wait for 20 ns;
			 X <="11010001";
			 wait for 20 ns;
			 X <="11010010";
			 wait for 20 ns;
			 X <="11010011";
			 wait for 20 ns;
			 X <="11010100";
			 wait for 20 ns;
			 X <="11010101";
			 wait for 20 ns;
			 X <="11010110";
			 wait for 20 ns;
			 X <="11010111";
			 wait for 20 ns;
			 X <="11011000";
			 wait for 20 ns;
			 X <="11011001";
			 wait for 20 ns;
			 X <="11011010";
			 wait for 20 ns;
			 X <="11011011";
			 wait for 20 ns;
			 X <="11011100";
			 wait for 20 ns;
			 X <="11011101";
			 wait for 20 ns;
			 X <="11011110";
			 wait for 20 ns;
			 X <="11011111";
			 wait for 20 ns;
			 X <="11100000";
			 wait for 20 ns;
			 X <="11100001";
			 wait for 20 ns;
			 X <="11100010";
			 wait for 20 ns;
			 X <="11100011";
			 wait for 20 ns;
			 X <="11100100";
			 wait for 20 ns;
			 X <="11100101";
			 wait for 20 ns;
			 X <="11100110";
			 wait for 20 ns;
			 X <="11100111";
			 wait for 20 ns;
			 X <="11101000";
			 wait for 20 ns;
			 X <="11101001";
			 wait for 20 ns;
			 X <="11101010";
			 wait for 20 ns;
			 X <="11101011";
			 wait for 20 ns;
			 X <="11101100";
			 wait for 20 ns;
			 X <="11101101";
			 wait for 20 ns;
			 X <="11101110";
			 wait for 20 ns;
			 X <="11101111";
			 wait for 20 ns;
			 X <="11110000";
			 wait for 20 ns;
			 X <="11110001";
			 wait for 20 ns;
			 X <="11110010";
			 wait for 20 ns;
			 X <="11110011";
			 wait for 20 ns;
			 X <="11110100";
			 wait for 20 ns;
			 X <="11110101";
			 wait for 20 ns;
			 X <="11110110";
			 wait for 20 ns;
			 X <="11110111";
			 wait for 20 ns;
			 X <="11111000";
			 wait for 20 ns;
			 X <="11111001";
			 wait for 20 ns;
			 X <="11111010";
			 wait for 20 ns;
			 X <="11111011";
			 wait for 20 ns;
			 X <="11111100";
			 wait for 20 ns;
			 X <="11111101";
			 wait for 20 ns;
			 X <="11111110";
			 wait for 20 ns;
			 X <="11111111";
			 wait for 20 ns;
	 end process; 
END SIMULATION; 
