-- Tabla de consulta de Datos
-- 
-- Diseño Lógico
-- Gustavo David Mendoza Pinto

LIBRARY IEEE; 
USE IEEE.std_logic_1164.all; 
Entity LUT_SIN_7SEG is 
	 port(
		 X : in  std_logic_vector(9 downto 0);
		 Y : out std_logic_vector(41 downto 0));
END LUT_SIN_7SEG; 
Architecture TABLE of LUT_SIN_7SEG is 
BEGIN 
	 process(X) 
	 begin 
		 case X is 
			 when "0000000000" => Y <= "000000011111101111110111111011111101111110"; -- Argumento 0( 0.0 Radianes) Función 0.0
			 when "0000000001" => Y <= "000000011111101111110111111000111110110000"; -- Argumento 1( 0.006135923151542565 Radianes) Función 0.006135884649154475
			 when "0000000010" => Y <= "000000011111101111110011000010011011001101"; -- Argumento 2( 0.01227184630308513 Radianes) Función 0.012271538285719925
			 when "0000000011" => Y <= "000000011111101111110011000011111110110011"; -- Argumento 3( 0.018407769454627694 Radianes) Función 0.01840672990580482
			 when "0000000100" => Y <= "000000011111101111110100110101100111011011"; -- Argumento 4( 0.02454369260617026 Radianes) Función 0.024541228522912288
			 when "0000000101" => Y <= "000000011111101111110111100111111100011111"; -- Argumento 5( 0.030679615757712823 Radianes) Función 0.030674803176636626
			 when "0000000110" => Y <= "000000011111101111110111100100111111111111"; -- Argumento 6( 0.03681553890925539 Radianes) Función 0.03680722294135883
			 when "0000000111" => Y <= "000000011111101111110011001110011011110011"; -- Argumento 7( 0.04295146206079795 Radianes) Función 0.04293825693494082
			 when "0000001000" => Y <= "000000011111101111110011001111100111111110"; -- Argumento 8( 0.04908738521234052 Radianes) Función 0.049067674327418015
			 when "0000001001" => Y <= "000000011111101111110101101110110110110000"; -- Argumento 9( 0.05522330836388308 Radianes) Función 0.05519524434968994
			 when "0000001010" => Y <= "000000011111101111110001111101100001111001"; -- Argumento 10( 0.06135923151542565 Radianes) Función 0.06132073630220858
			 when "0000001011" => Y <= "000000011111101111110001111111100010110011"; -- Argumento 11( 0.0674951546669682 Radianes) Función 0.06744391956366405
			 when "0000001100" => Y <= "000000011111101111110111000111110011011011"; -- Argumento 12( 0.07363107781851078 Radianes) Función 0.07356456359966743
			 when "0000001101" => Y <= "000000011111101111110111000111100110011111"; -- Argumento 13( 0.07976700097005335 Radianes) Función 0.07968243797143013
			 when "0000001110" => Y <= "000000011111101111110111111110110111110001"; -- Argumento 14( 0.0859029241215959 Radianes) Función 0.0857973123444399
			 when "0000001111" => Y <= "000000011111101111110111001101100001110011"; -- Argumento 15( 0.09203884727313846 Radianes) Función 0.09190895649713272
			 when "0000010000" => Y <= "000000011111101111110111001111111111111110"; -- Argumento 16( 0.09817477042468103 Radianes) Función 0.0980171403295606
			 when "0000010001" => Y <= "000000011111100110000111111001100110110000"; -- Argumento 17( 0.1043106935762236 Radianes) Función 0.10412163387205459
			 when "0000010010" => Y <= "000000011111100110000011000011111101001101"; -- Argumento 18( 0.11044661672776616 Radianes) Función 0.11022220729388306
			 when "0000010011" => Y <= "000000011111100110000011000000111111111001"; -- Argumento 19( 0.11658253987930872 Radianes) Función 0.11631863091190475
			 when "0000010100" => Y <= "000000011111100110000100110110011010110011"; -- Argumento 20( 0.1227184630308513 Radianes) Función 0.1224106751992162
			 when "0000010101" => Y <= "000000011111100110000100110111111110110011"; -- Argumento 21( 0.12885438618239387 Radianes) Función 0.12849811079379317
			 when "0000010110" => Y <= "000000011111100110000111100101100111011011"; -- Argumento 22( 0.1349903093339364 Radianes) Función 0.13458070850712617
			 when "0000010111" => Y <= "000000011111100110000011001111111100011111"; -- Argumento 23( 0.14112623248547898 Radianes) Función 0.1406582393328492
			 when "0000011000" => Y <= "000000011111100110000011001100111111110001"; -- Argumento 24( 0.14726215563702155 Radianes) Función 0.14673047445536175
			 when "0000011001" => Y <= "000000011111100110000101101110011011110001"; -- Argumento 25( 0.15339807878856412 Radianes) Función 0.15279718525844344
			 when "0000011010" => Y <= "000000011111100110000101101111111111111111"; -- Argumento 26( 0.1595340019401067 Radianes) Función 0.15885814333386145
			 when "0000011011" => Y <= "000000011111100110000001111101100111110011"; -- Argumento 27( 0.16566992509164924 Radianes) Función 0.16491312048996992
			 when "0000011100" => Y <= "000000011111100110000111000111111101110011"; -- Argumento 28( 0.1718058482431918 Radianes) Función 0.17096188876030122
			 when "0000011101" => Y <= "000000011111100110000111000111100011111110"; -- Argumento 29( 0.17794177139473438 Radianes) Función 0.17700422041214875
			 when "0000011110" => Y <= "000000011111100110000111111111110011111110"; -- Argumento 30( 0.18407769454627693 Radianes) Función 0.18303988795514095
			 when "0000011111" => Y <= "000000011111100110000111111111100111111110"; -- Argumento 31( 0.1902136176978195 Radianes) Función 0.1890686641498062
			 when "0000100000" => Y <= "000000011111100110000111001110110111111110"; -- Argumento 32( 0.19634954084936207 Radianes) Función 0.19509032201612825
			 when "0000100001" => Y <= "000000011111101001101111111001100000110000"; -- Argumento 33( 0.20248546400090464 Radianes) Función 0.2011046348420919
			 when "0000100010" => Y <= "000000011111101001101111111011100010110000"; -- Argumento 34( 0.2086213871524472 Radianes) Función 0.20711137619221856
			 when "0000100011" => Y <= "000000011111101001101011000011110010110000"; -- Argumento 35( 0.21475731030398976 Radianes) Función 0.21311031991609136
			 when "0000100100" => Y <= "000000011111101001101011000011100110110000"; -- Argumento 36( 0.22089323345553233 Radianes) Función 0.2191012401568698
			 when "0000100101" => Y <= "000000011111101001101100110110110111111110"; -- Argumento 37( 0.2270291566070749 Radianes) Función 0.22508391135979283
			 when "0000100110" => Y <= "000000011111101001101111100101100001111110"; -- Argumento 38( 0.23316507975861744 Radianes) Función 0.2310581082806711
			 when "0000100111" => Y <= "000000011111101001101111100111100011111110"; -- Argumento 39( 0.23930100291016002 Radianes) Función 0.2370236059943672
			 when "0000101000" => Y <= "000000011111101001101011001110011011110011"; -- Argumento 40( 0.2454369260617026 Radianes) Función 0.24298017990326387
			 when "0000101001" => Y <= "000000011111101001101011001111111111110011"; -- Argumento 41( 0.25157284921324513 Radianes) Función 0.24892760574572015
			 when "0000101010" => Y <= "000000011111101001101101101101100111111111"; -- Argumento 42( 0.25770877236478773 Radianes) Función 0.25486565960451457
			 when "0000101011" => Y <= "000000011111101001101001111111111101110001"; -- Argumento 43( 0.2638446955163303 Radianes) Función 0.2607941179152755
			 when "0000101100" => Y <= "000000011111101001101001111100111111110001"; -- Argumento 44( 0.2699806186678728 Radianes) Función 0.26671275747489837
			 when "0000101101" => Y <= "000000011111101001101111000110011010011111"; -- Argumento 45( 0.2761165418194154 Radianes) Función 0.272621355449949
			 when "0000101110" => Y <= "000000011111101001101111000111111111011011"; -- Argumento 46( 0.28225246497095796 Radianes) Función 0.27851968938505306
			 when "0000101111" => Y <= "000000011111101001101111111101100110110011"; -- Argumento 47( 0.28838838812250056 Radianes) Función 0.2844075372112719
			 when "0000110000" => Y <= "000000011111101001101111001111111101001101"; -- Argumento 48( 0.2945243112740431 Radianes) Función 0.29028467725446233
			 when "0000110001" => Y <= "000000011111101001101111001100111110110000"; -- Argumento 49( 0.30066023442558565 Radianes) Función 0.2961508882436238
			 when "0000110010" => Y <= "000000011111101111001111111010011011111110"; -- Argumento 50( 0.30679615757712825 Radianes) Función 0.3020059493192281
			 when "0000110011" => Y <= "000000011111101111001111111011100011111111"; -- Argumento 51( 0.3129320807286708 Radianes) Función 0.30784964004153487
			 when "0000110100" => Y <= "000000011111101111001011000011110010011111"; -- Argumento 52( 0.3190680038802134 Radianes) Función 0.3136817403988915
			 when "0000110101" => Y <= "000000011111101111001011000011100111011011"; -- Argumento 53( 0.32520392703175593 Radianes) Función 0.3195020308160157
			 when "0000110110" => Y <= "000000011111101111001100110110110111111001"; -- Argumento 54( 0.3313398501832985 Radianes) Función 0.3253102921622629
			 when "0000110111" => Y <= "000000011111101111001111100101100000110000"; -- Argumento 55( 0.3374757733348411 Radianes) Función 0.33110630575987643
			 when "0000111000" => Y <= "000000011111101111001111100100111111111111"; -- Argumento 56( 0.3436116964863836 Radianes) Función 0.33688985339222005
			 when "0000111001" => Y <= "000000011111101111001011001110011010011111"; -- Argumento 57( 0.34974761963792617 Radianes) Función 0.3426607173119944
			 when "0000111010" => Y <= "000000011111101111001011001111111110110011"; -- Argumento 58( 0.35588354278946877 Radianes) Función 0.34841868024943456
			 when "0000111011" => Y <= "000000011111101111001101101101100110110000"; -- Argumento 59( 0.3620194659410113 Radianes) Función 0.35416352542049034
			 when "0000111100" => Y <= "000000011111101111001101101111100111111111"; -- Argumento 60( 0.36815538909255385 Radianes) Función 0.3598950365349881
			 when "0000111101" => Y <= "000000011111101111001001111110110110011111"; -- Argumento 61( 0.37429131224409645 Radianes) Función 0.36561299780477385
			 when "0000111110" => Y <= "000000011111101111001111000101100001111001"; -- Argumento 62( 0.380427235395639 Radianes) Función 0.37131719395183754
			 when "0000111111" => Y <= "000000011111101111001111000111100011111110"; -- Argumento 63( 0.3865631585471816 Radianes) Función 0.37700741021641826
			 when "0001000000" => Y <= "000000011111101111001111111110011010011111"; -- Argumento 64( 0.39269908169872414 Radianes) Función 0.3826834323650898
			 when "0001000001" => Y <= "000000011111101111001111111111111111111001"; -- Argumento 65( 0.3988350048502667 Radianes) Función 0.38834504669882625
			 when "0001000010" => Y <= "000000011111101111001111001111110011110011"; -- Argumento 66( 0.4049709280018093 Radianes) Función 0.3939920400610481
			 when "0001000011" => Y <= "000000011111101111001111001111100110011111"; -- Argumento 67( 0.4111068511533518 Radianes) Función 0.3996241998456468
			 when "0001000100" => Y <= "000000011111100110011111111010110111001101"; -- Argumento 68( 0.4172427743048944 Radianes) Función 0.40524131400498986
			 when "0001000101" => Y <= "000000011111100110011011000011111101111111"; -- Argumento 69( 0.42337869745643697 Radianes) Función 0.4108431710579039
			 when "0001000110" => Y <= "000000011111100110011011000000111110110011"; -- Argumento 70( 0.4295146206079795 Radianes) Función 0.41642956009763715
			 when "0001000111" => Y <= "000000011111100110011100110110011011111110"; -- Argumento 71( 0.4356505437595221 Radianes) Función 0.4220002707997997
			 when "0001001000" => Y <= "000000011111100110011100110111100011011011"; -- Argumento 72( 0.44178646691106466 Radianes) Función 0.4275550934302821
			 when "0001001001" => Y <= "000000011111100110011111100111110011111110"; -- Argumento 73( 0.4479223900626072 Radianes) Función 0.43309381885315196
			 when "0001001010" => Y <= "000000011111100110011111100111111110011111"; -- Argumento 74( 0.4540583132141498 Radianes) Función 0.43861623853852766
			 when "0001001011" => Y <= "000000011111100110011011001101100110110000"; -- Argumento 75( 0.46019423636569234 Radianes) Función 0.4441221445704292
			 when "0001001100" => Y <= "000000011111100110011011001111100110011111"; -- Argumento 76( 0.4663301595172349 Radianes) Función 0.44961132965460654
			 when "0001001101" => Y <= "000000011111100110011101101110110111111110"; -- Argumento 77( 0.4724660826687775 Radianes) Función 0.45508358712634384
			 when "0001001110" => Y <= "000000011111100110011001111111111101011011"; -- Argumento 78( 0.47860200582032003 Radianes) Función 0.46053871095824
			 when "0001001111" => Y <= "000000011111100110011001111110110111110011"; -- Argumento 79( 0.48473792897186263 Radianes) Función 0.4659764957679662
			 when "0001010000" => Y <= "000000011111100110011111000101100001111001"; -- Argumento 80( 0.4908738521234052 Radianes) Función 0.47139673682599764
			 when "0001010001" => Y <= "000000011111100110011111000100111111110001"; -- Argumento 81( 0.4970097752749477 Radianes) Función 0.4767992300633221
			 when "0001010010" => Y <= "000000011111100110011111111110011010110000"; -- Argumento 82( 0.5031456984264903 Radianes) Función 0.4821837720791227
			 when "0001010011" => Y <= "000000011111100110011111111111100011011011"; -- Argumento 83( 0.5092816215780329 Radianes) Función 0.487550160148436
			 when "0001010100" => Y <= "000000011111100110011111001110011011111111"; -- Argumento 84( 0.5154175447295755 Radianes) Función 0.49289819222978404
			 when "0001010101" => Y <= "000000011111100110011111001111111111001101"; -- Argumento 85( 0.521553467881118 Radianes) Función 0.49822766697278187
			 when "0001010110" => Y <= "000000011111101011011111111011110011011011"; -- Argumento 86( 0.5276893910326605 Radianes) Función 0.5035383837257176
			 when "0001010111" => Y <= "000000011111101011011111111011111111111111"; -- Argumento 87( 0.5338253141842031 Radianes) Función 0.508830142543107
			 when "0001011000" => Y <= "000000011111101011011011000001100110110000"; -- Argumento 88( 0.5399612373357456 Radianes) Función 0.5141027441932217
			 when "0001011001" => Y <= "000000011111101011011011000011100111111001"; -- Argumento 89( 0.5460971604872883 Radianes) Función 0.5193559901655896
			 when "0001011010" => Y <= "000000011111101011011100110101100111011011"; -- Argumento 90( 0.5522330836388308 Radianes) Función 0.524589682678469
			 when "0001011011" => Y <= "000000011111101011011100110111100111111111"; -- Argumento 91( 0.5583690067903734 Radianes) Función 0.5298036246862946
			 when "0001011100" => Y <= "000000011111101011011111100101100111110011"; -- Argumento 92( 0.5645049299419159 Radianes) Función 0.5349976198870972
			 when "0001011101" => Y <= "000000011111101011011011001111111100110000"; -- Argumento 93( 0.5706408530934585 Radianes) Función 0.5401714727298929
			 when "0001011110" => Y <= "000000011111101011011011001110110111111001"; -- Argumento 94( 0.5767767762450011 Radianes) Función 0.5453249884220465
			 when "0001011111" => Y <= "000000011111101011011101101111111100110011"; -- Argumento 95( 0.5829126993965437 Radianes) Función 0.5504579729366048
			 when "0001100000" => Y <= "000000011111101011011101101110110111011011"; -- Argumento 96( 0.5890486225480862 Radianes) Función 0.5555702330196022
			 when "0001100001" => Y <= "000000011111101011011001111111111100011111"; -- Argumento 97( 0.5951845456996288 Radianes) Función 0.560661576197336
			 when "0001100010" => Y <= "000000011111101011011001111110110111110001"; -- Argumento 98( 0.6013204688511713 Radianes) Función 0.5657318107836131
			 when "0001100011" => Y <= "000000011111101011011111000111111101110001"; -- Argumento 99( 0.607456392002714 Radianes) Función 0.5707807458869673
			 when "0001100100" => Y <= "000000011111101011011111000110110111111111"; -- Argumento 100( 0.6135923151542565 Radianes) Función 0.5758081914178453
			 when "0001100101" => Y <= "000000011111101011011111111111111101111111"; -- Argumento 101( 0.619728238305799 Radianes) Función 0.5808139580957645
			 when "0001100110" => Y <= "000000011111101011011111111110110111110001"; -- Argumento 102( 0.6258641614573416 Radianes) Función 0.5857978574564389
			 when "0001100111" => Y <= "000000011111101011011111001111111101110001"; -- Argumento 103( 0.6320000846088841 Radianes) Función 0.5907597018588742
			 when "0001101000" => Y <= "000000011111101011011111001110110110011111"; -- Argumento 104( 0.6381360077604268 Radianes) Función 0.5956993044924334
			 when "0001101001" => Y <= "000000011111100011111111111011111100011111"; -- Argumento 105( 0.6442719309119693 Radianes) Función 0.600616479383869
			 when "0001101010" => Y <= "000000011111100011111111111010110111011011"; -- Argumento 106( 0.6504078540635119 Radianes) Función 0.6055110414043255
			 when "0001101011" => Y <= "000000011111100011111011000011111101111001"; -- Argumento 107( 0.6565437772150544 Radianes) Función 0.6103828062763095
			 when "0001101100" => Y <= "000000011111100011111011000010110111001101"; -- Argumento 108( 0.662679700366597 Radianes) Función 0.6152315905806268
			 when "0001101101" => Y <= "000000011111100011111100110111111101111110"; -- Argumento 109( 0.6688156235181395 Radianes) Función 0.6200572117632891
			 when "0001101110" => Y <= "000000011111100011111100110101100111111111"; -- Argumento 110( 0.6749515466696822 Radianes) Función 0.6248594881423863
			 when "0001101111" => Y <= "000000011111100011111100110111100110011111"; -- Argumento 111( 0.6810874698212247 Radianes) Función 0.629638238914927
			 when "0001110000" => Y <= "000000011111100011111111100101100111111001"; -- Argumento 112( 0.6872233929727672 Radianes) Función 0.6343932841636455
			 when "0001110001" => Y <= "000000011111100011111111100111100110110000"; -- Argumento 113( 0.6933593161243098 Radianes) Función 0.6391244448637757
			 when "0001110010" => Y <= "000000011111100011111011001111110011111111"; -- Argumento 114( 0.6994952392758523 Radianes) Función 0.6438315428897914
			 when "0001110011" => Y <= "000000011111100011111011001111111111011011"; -- Argumento 115( 0.705631162427395 Radianes) Función 0.6485144010221124
			 when "0001110100" => Y <= "000000011111100011111101101111110010110000"; -- Argumento 116( 0.7117670855789375 Radianes) Función 0.6531728429537768
			 when "0001110101" => Y <= "000000011111100011111101101111100011111111"; -- Argumento 117( 0.7179030087304801 Radianes) Función 0.6578066932970786
			 when "0001110110" => Y <= "000000011111100011111001111110011010110011"; -- Argumento 118( 0.7240389318820226 Radianes) Función 0.6624157775901718
			 when "0001110111" => Y <= "000000011111100011111001111100111111110011"; -- Argumento 119( 0.7301748550335652 Radianes) Función 0.6669999223036375
			 when "0001111000" => Y <= "000000011111100011111111000101100001011011"; -- Argumento 120( 0.7363107781851077 Radianes) Función 0.6715589548470183
			 when "0001111001" => Y <= "000000011111100011111111000100111111111110"; -- Argumento 121( 0.7424467013366504 Radianes) Función 0.6760927035753159
			 when "0001111010" => Y <= "000000011111100011111111111111111100011111"; -- Argumento 122( 0.7485826244881929 Radianes) Función 0.680600997795453
			 when "0001111011" => Y <= "000000011111100011111111111110110111111110"; -- Argumento 123( 0.7547185476397354 Radianes) Función 0.6850836677727004
			 when "0001111100" => Y <= "000000011111100011111111111111100111011011"; -- Argumento 124( 0.760854470791278 Radianes) Función 0.6895405447370669
			 when "0001111101" => Y <= "000000011111100011111111001111110011110011"; -- Argumento 125( 0.7669903939428205 Radianes) Función 0.693971460889654
			 when "0001111110" => Y <= "000000011111100011111111001111111111111001"; -- Argumento 126( 0.7731263170943632 Radianes) Función 0.6983762494089729
			 when "0001111111" => Y <= "000000011111101110001111111010011011110001"; -- Argumento 127( 0.7792622402459057 Radianes) Función 0.7027547444572253
			 when "0010000000" => Y <= "000000011111101110001111111011100010110000"; -- Argumento 128( 0.7853981633974483 Radianes) Función 0.7071067811865475
			 when "0010000001" => Y <= "000000011111101110001011000001100000110011"; -- Argumento 129( 0.7915340865489908 Radianes) Función 0.7114321957452164
			 when "0010000010" => Y <= "000000011111101110001011000010110111110001"; -- Argumento 130( 0.7976700097005334 Radianes) Función 0.7157308252838186
			 when "0010000011" => Y <= "000000011111101110001100110111111101111110"; -- Argumento 131( 0.803805932852076 Radianes) Función 0.7200025079613817
			 when "0010000100" => Y <= "000000011111101110001100110101100111001101"; -- Argumento 132( 0.8099418560036186 Radianes) Función 0.7242470829514669
			 when "0010000101" => Y <= "000000011111101110001100110111111110110011"; -- Argumento 133( 0.8160777791551611 Radianes) Función 0.7284643904482252
			 when "0010000110" => Y <= "000000011111101110001111100110011010011111"; -- Argumento 134( 0.8222137023067037 Radianes) Función 0.7326542716724128
			 when "0010000111" => Y <= "000000011111101110001111100100111111111111"; -- Argumento 135( 0.8283496254582462 Radianes) Función 0.7368165688773698
			 when "0010001000" => Y <= "000000011111101110001011001111111101110011"; -- Argumento 136( 0.8344855486097889 Radianes) Función 0.7409511253549591
			 when "0010001001" => Y <= "000000011111101110001011001110110111111110"; -- Argumento 137( 0.8406214717613314 Radianes) Función 0.745057785441466
			 when "0010001010" => Y <= "000000011111101110001011001111100110110000"; -- Argumento 138( 0.8467573949128739 Radianes) Función 0.7491363945234593
			 when "0010001011" => Y <= "000000011111101110001101101111110010110000"; -- Argumento 139( 0.8528933180644165 Radianes) Función 0.7531867990436124
			 when "0010001100" => Y <= "000000011111101110001101101111100011001101"; -- Argumento 140( 0.859029241215959 Radianes) Función 0.7572088465064845
			 when "0010001101" => Y <= "000000011111101110001001111101100001001101"; -- Argumento 141( 0.8651651643675016 Radianes) Función 0.7612023854842617
			 when "0010001110" => Y <= "000000011111101110001001111110110110110000"; -- Argumento 142( 0.8713010875190442 Radianes) Función 0.765167265622459
			 when "0010001111" => Y <= "000000011111101110001001111111100110110000"; -- Argumento 143( 0.8774370106705868 Radianes) Función 0.7691033376455796
			 when "0010010000" => Y <= "000000011111101110001111000111110011111110"; -- Argumento 144( 0.8835729338221293 Radianes) Función 0.7730104533627369
			 when "0010010001" => Y <= "000000011111101110001111000100111111111111"; -- Argumento 145( 0.8897088569736719 Radianes) Función 0.7768884656732323
			 when "0010010010" => Y <= "000000011111101110001111111111111101110001"; -- Argumento 146( 0.8958447801252144 Radianes) Función 0.7807372285720944
			 when "0010010011" => Y <= "000000011111101110001111111101100111011011"; -- Argumento 147( 0.9019807032767571 Radianes) Función 0.7845565971555752
			 when "0010010100" => Y <= "000000011111101110001111111111111111111001"; -- Argumento 148( 0.9081166264282996 Radianes) Función 0.7883464276266062
			 when "0010010101" => Y <= "000000011111101110001111001110011010110000"; -- Argumento 149( 0.9142525495798421 Radianes) Función 0.7921065773002123
			 when "0010010110" => Y <= "000000011111101110001111001110110111111111"; -- Argumento 150( 0.9203884727313847 Radianes) Función 0.7958369046088835
			 when "0010010111" => Y <= "000000011111101110001111001111100111011011"; -- Argumento 151( 0.9265243958829272 Radianes) Función 0.7995372691079049
			 when "0010011000" => Y <= "000000011111101111111111111011110011001101"; -- Argumento 152( 0.9326603190344698 Radianes) Función 0.8032075314806448
			 when "0010011001" => Y <= "000000011111101111111111111000111111111111"; -- Argumento 153( 0.9387962421860124 Radianes) Función 0.8068475535437992
			 when "0010011010" => Y <= "000000011111101111111011000011111100110011"; -- Argumento 154( 0.944932165337555 Radianes) Función 0.8104571982525948
			 when "0010011011" => Y <= "000000011111101111111011000001100111111110"; -- Argumento 155( 0.9510680884890975 Radianes) Función 0.8140363297059483
			 when "0010011100" => Y <= "000000011111101111111011000011100011011011"; -- Argumento 156( 0.9572040116406401 Radianes) Función 0.8175848131515836
			 when "0010011101" => Y <= "000000011111101111111100110101100000110000"; -- Argumento 157( 0.9633399347921826 Radianes) Función 0.8211025149911046
			 when "0010011110" => Y <= "000000011111101111111100110101100111011011"; -- Argumento 158( 0.9694758579437253 Radianes) Función 0.8245893027850253
			 when "0010011111" => Y <= "000000011111101111111100110111111111111110"; -- Argumento 159( 0.9756117810952678 Radianes) Función 0.8280450452577557
			 when "0010100000" => Y <= "000000011111101111111111100101100000110011"; -- Argumento 160( 0.9817477042468103 Radianes) Función 0.8314696123025452
			 when "0010100001" => Y <= "000000011111101111111111100101100111111111"; -- Argumento 161( 0.9878836273983529 Radianes) Función 0.83486287498638
			 when "0010100010" => Y <= "000000011111101111111111100111111111001101"; -- Argumento 162( 0.9940195505498954 Radianes) Función 0.838224705554838
			 when "0010100011" => Y <= "000000011111101111111011001101100001011011"; -- Argumento 163( 1.000155473701438 Radianes) Función 0.8415549774368983
			 when "0010100100" => Y <= "000000011111101111111011001101100111111111"; -- Argumento 164( 1.0062913968529805 Radianes) Función 0.844853565249707
			 when "0010100101" => Y <= "000000011111101111111011001111111110110000"; -- Argumento 165( 1.012427320004523 Radianes) Función 0.8481203448032971
			 when "0010100110" => Y <= "000000011111101111111101101101100001111001"; -- Argumento 166( 1.0185632431560658 Radianes) Función 0.8513551931052652
			 when "0010100111" => Y <= "000000011111101111111101101101100111011011"; -- Argumento 167( 1.0246991663076084 Radianes) Función 0.8545579883654005
			 when "0010101000" => Y <= "000000011111101111111101101111100011110001"; -- Argumento 168( 1.030835089459151 Radianes) Función 0.857728610000272
			 when "0010101001" => Y <= "000000011111101111111001111111111101111111"; -- Argumento 169( 1.0369710126106935 Radianes) Función 0.8608669386377672
			 when "0010101010" => Y <= "000000011111101111111001111111110011110011"; -- Argumento 170( 1.043106935762236 Radianes) Función 0.8639728561215867
			 when "0010101011" => Y <= "000000011111101111111001111111100011111110"; -- Argumento 171( 1.0492428589137786 Radianes) Función 0.8670462455156925
			 when "0010101100" => Y <= "000000011111101111111111000111111101111110"; -- Argumento 172( 1.055378782065321 Radianes) Función 0.8700869911087113
			 when "0010101101" => Y <= "000000011111101111111111000111110011111110"; -- Argumento 173( 1.0615147052168636 Radianes) Función 0.87309497841829
			 when "0010101110" => Y <= "000000011111101111111111000100111111111110"; -- Argumento 174( 1.0676506283684062 Radianes) Función 0.8760700941954065
			 when "0010101111" => Y <= "000000011111101111111111000111100111111110"; -- Argumento 175( 1.0737865515199487 Radianes) Función 0.8790122264286334
			 when "0010110000" => Y <= "000000011111101111111111111101100001110011"; -- Argumento 176( 1.0799224746714913 Radianes) Función 0.8819212643483549
			 when "0010110001" => Y <= "000000011111101111111111111101100111110001"; -- Argumento 177( 1.086058397823034 Radianes) Función 0.8847970984309378
			 when "0010110010" => Y <= "000000011111101111111111111111100010011111"; -- Argumento 178( 1.0921943209745766 Radianes) Función 0.8876396204028539
			 when "0010110011" => Y <= "000000011111101111111111001111111100110011"; -- Argumento 179( 1.0983302441261191 Radianes) Función 0.8904487232447579
			 when "0010110100" => Y <= "000000011111101111111111001111110011001101"; -- Argumento 180( 1.1044661672776617 Radianes) Función 0.8932243011955153
			 when "0010110101" => Y <= "000000011111101111111111001110110111110011"; -- Argumento 181( 1.1106020904292042 Radianes) Función 0.8959662497561851
			 when "0010110110" => Y <= "000000011111101111111111001111111110011111"; -- Argumento 182( 1.1167380135807468 Radianes) Función 0.8986744656939538
			 when "0010110111" => Y <= "000000011111101110011111111001100001111001"; -- Argumento 183( 1.1228739367322893 Radianes) Función 0.901348847046022
			 when "0010111000" => Y <= "000000011111101110011111111011110011110011"; -- Argumento 184( 1.1290098598838318 Radianes) Función 0.9039892931234433
			 when "0010111001" => Y <= "000000011111101110011111111000111111011011"; -- Argumento 185( 1.1351457830353744 Radianes) Función 0.9065957045149153
			 when "0010111010" => Y <= "000000011111101110011111111011100110110000"; -- Argumento 186( 1.141281706186917 Radianes) Función 0.9091679830905224
			 when "0010111011" => Y <= "000000011111101110011011000001100001110001"; -- Argumento 187( 1.1474176293384597 Radianes) Función 0.9117060320054299
			 when "0010111100" => Y <= "000000011111101110011011000001100111001101"; -- Argumento 188( 1.1535535524900022 Radianes) Función 0.9142097557035307
			 when "0010111101" => Y <= "000000011111101110011011000000111110011111"; -- Argumento 189( 1.1596894756415448 Radianes) Función 0.9166790599210427
			 when "0010111110" => Y <= "000000011111101110011011000011100110110000"; -- Argumento 190( 1.1658253987930873 Radianes) Función 0.9191138516900578
			 when "0010111111" => Y <= "000000011111101110011100110101100001011011"; -- Argumento 191( 1.1719613219446299 Radianes) Función 0.9215140393420419
			 when "0011000000" => Y <= "000000011111101110011100110111110011111111"; -- Argumento 192( 1.1780972450961724 Radianes) Función 0.9238795325112867
			 when "0011000001" => Y <= "000000011111101110011100110100111111001101"; -- Argumento 193( 1.184233168247715 Radianes) Función 0.9262102421383114
			 when "0011000010" => Y <= "000000011111101110011100110111111111011011"; -- Argumento 194( 1.1903690913992575 Radianes) Función 0.9285060804732156
			 when "0011000011" => Y <= "000000011111101110011111100111111101110001"; -- Argumento 195( 1.1965050145508 Radianes) Función 0.9307669610789837
			 when "0011000100" => Y <= "000000011111101110011111100110011011110011"; -- Argumento 196( 1.2026409377023426 Radianes) Función 0.9329927988347388
			 when "0011000101" => Y <= "000000011111101110011111100110110110110000"; -- Argumento 197( 1.2087768608538851 Radianes) Función 0.9351835099389475
			 when "0011000110" => Y <= "000000011111101110011111100111100011111001"; -- Argumento 198( 1.214912784005428 Radianes) Función 0.937339011912575
			 when "0011000111" => Y <= "000000011111101110011111100111100110110011"; -- Argumento 199( 1.2210487071569704 Radianes) Función 0.9394592236021899
			 when "0011001000" => Y <= "000000011111101110011011001101100001011011"; -- Argumento 200( 1.227184630308513 Radianes) Función 0.9415440651830208
			 when "0011001001" => Y <= "000000011111101110011011001111110011011011"; -- Argumento 201( 1.2333205534600555 Radianes) Función 0.9435934581619604
			 when "0011001010" => Y <= "000000011111101110011011001110110110011111"; -- Argumento 202( 1.239456476611598 Radianes) Función 0.9456073253805213
			 when "0011001011" => Y <= "000000011111101110011011001111100011011011"; -- Argumento 203( 1.2455923997631406 Radianes) Función 0.9475855910177411
			 when "0011001100" => Y <= "000000011111101110011011001111100111011011"; -- Argumento 204( 1.2517283229146832 Radianes) Función 0.9495281805930367
			 when "0011001101" => Y <= "000000011111101110011101101101100000110011"; -- Argumento 205( 1.2578642460662257 Radianes) Función 0.9514350209690083
			 when "0011001110" => Y <= "000000011111101110011101101111110011111001"; -- Argumento 206( 1.2640001692177683 Radianes) Función 0.9533060403541938
			 when "0011001111" => Y <= "000000011111101110011101101110110110110000"; -- Argumento 207( 1.2701360923693108 Radianes) Función 0.9551411683057707
			 when "0011010000" => Y <= "000000011111101110011101101100111111110011"; -- Argumento 208( 1.2762720155208536 Radianes) Función 0.9569403357322089
			 when "0011010001" => Y <= "000000011111101110011101101111111111110001"; -- Argumento 209( 1.282407938672396 Radianes) Función 0.9587034748958716
			 when "0011010010" => Y <= "000000011111101110011001111111111100110011"; -- Argumento 210( 1.2885438618239387 Radianes) Función 0.9604305194155658
			 when "0011010011" => Y <= "000000011111101110011001111110011010110000"; -- Argumento 211( 1.2946797849754812 Radianes) Función 0.9621214042690416
			 when "0011010100" => Y <= "000000011111101110011001111111110011110001"; -- Argumento 212( 1.3008157081270237 Radianes) Función 0.9637760657954398
			 when "0011010101" => Y <= "000000011111101110011001111110110111111001"; -- Argumento 213( 1.3069516312785663 Radianes) Función 0.9653944416976894
			 when "0011010110" => Y <= "000000011111101110011001111100111111110011"; -- Argumento 214( 1.3130875544301088 Radianes) Función 0.9669764710448521
			 when "0011010111" => Y <= "000000011111101110011001111111111111011011"; -- Argumento 215( 1.3192234775816514 Radianes) Función 0.9685220942744173
			 when "0011011000" => Y <= "000000011111101110011111000111111101111110"; -- Argumento 216( 1.325359400733194 Radianes) Función 0.970031253194544
			 when "0011011001" => Y <= "000000011111101110011111000101100001011011"; -- Argumento 217( 1.3314953238847365 Radianes) Función 0.9715038909862518
			 when "0011011010" => Y <= "000000011111101110011111000110011011110011"; -- Argumento 218( 1.337631247036279 Radianes) Función 0.9729399522055601
			 when "0011011011" => Y <= "000000011111101110011111000101100111111001"; -- Argumento 219( 1.3437671701878218 Radianes) Función 0.9743393827855759
			 when "0011011100" => Y <= "000000011111101110011111000110110111110001"; -- Argumento 220( 1.3499030933393643 Radianes) Función 0.9757021300385286
			 when "0011011101" => Y <= "000000011111101110011111000111100011111110"; -- Argumento 221( 1.3560390164909069 Radianes) Función 0.9770281426577544
			 when "0011011110" => Y <= "000000011111101110011111000111111111111001"; -- Argumento 222( 1.3621749396424494 Radianes) Función 0.9783173707196277
			 when "0011011111" => Y <= "000000011111101110011111000111100111011011"; -- Argumento 223( 1.368310862793992 Radianes) Función 0.9795697656854405
			 when "0011100000" => Y <= "000000011111101110011111111111111101110001"; -- Argumento 224( 1.3744467859455345 Radianes) Función 0.9807852804032304
			 when "0011100001" => Y <= "000000011111101110011111111101100001110011"; -- Argumento 225( 1.380582709097077 Radianes) Función 0.9819638691095552
			 when "0011100010" => Y <= "000000011111101110011111111111110010110000"; -- Argumento 226( 1.3867186322486196 Radianes) Función 0.9831054874312163
			 when "0011100011" => Y <= "000000011111101110011111111101100111001101"; -- Argumento 227( 1.3928545554001621 Radianes) Función 0.984210092386929
			 when "0011100100" => Y <= "000000011111101110011111111110110111001101"; -- Argumento 228( 1.3989904785517047 Radianes) Función 0.9852776423889412
			 when "0011100101" => Y <= "000000011111101110011111111100111111111001"; -- Argumento 229( 1.4051264017032472 Radianes) Función 0.9863080972445987
			 when "0011100110" => Y <= "000000011111101110011111111111100011111001"; -- Argumento 230( 1.41126232485479 Radianes) Función 0.9873014181578584
			 when "0011100111" => Y <= "000000011111101110011111111111111111001101"; -- Argumento 231( 1.4173982480063325 Radianes) Función 0.9882575677307495
			 when "0011101000" => Y <= "000000011111101110011111111111100110110000"; -- Argumento 232( 1.423534171157875 Radianes) Función 0.989176509964781
			 when "0011101001" => Y <= "000000011111101110011111001111111101111110"; -- Argumento 233( 1.4296700943094176 Radianes) Función 0.9900582102622971
			 when "0011101010" => Y <= "000000011111101110011111001111111101110011"; -- Argumento 234( 1.4358060174609601 Radianes) Función 0.99090263542778
			 when "0011101011" => Y <= "000000011111101110011111001101100001110001"; -- Argumento 235( 1.4419419406125027 Radianes) Función 0.9917097536690995
			 when "0011101100" => Y <= "000000011111101110011111001110011010110011"; -- Argumento 236( 1.4480778637640452 Radianes) Función 0.99247953459871
			 when "0011101101" => Y <= "000000011111101110011111001111110011001101"; -- Argumento 237( 1.4542137869155878 Radianes) Función 0.9932119492347945
			 when "0011101110" => Y <= "000000011111101110011111001111110011110011"; -- Argumento 238( 1.4603497100671303 Radianes) Función 0.9939069700023561
			 when "0011101111" => Y <= "000000011111101110011111001101100111011011"; -- Argumento 239( 1.4664856332186729 Radianes) Función 0.9945645707342554
			 when "0011110000" => Y <= "000000011111101110011111001110110110110000"; -- Argumento 240( 1.4726215563702154 Radianes) Función 0.9951847266721968
			 when "0011110001" => Y <= "000000011111101110011111001110110111110001"; -- Argumento 241( 1.4787574795217582 Radianes) Función 0.9957674144676598
			 when "0011110010" => Y <= "000000011111101110011111001100111111111001"; -- Argumento 242( 1.4848934026733007 Radianes) Función 0.996312612182778
			 when "0011110011" => Y <= "000000011111101110011111001100111111111111"; -- Argumento 243( 1.4910293258248433 Radianes) Función 0.9968202992911657
			 when "0011110100" => Y <= "000000011111101110011111001111100011001101"; -- Argumento 244( 1.4971652489763858 Radianes) Función 0.9972904566786902
			 when "0011110101" => Y <= "000000011111101110011111001111100011110001"; -- Argumento 245( 1.5033011721279284 Radianes) Función 0.9977230666441916
			 when "0011110110" => Y <= "000000011111101110011111001111111110110000"; -- Argumento 246( 1.509437095279471 Radianes) Función 0.9981181129001492
			 when "0011110111" => Y <= "000000011111101110011111001111111110110011"; -- Argumento 247( 1.5155730184310134 Radianes) Función 0.9984755805732948
			 when "0011111000" => Y <= "000000011111101110011111001111111111110001"; -- Argumento 248( 1.521708941582556 Radianes) Función 0.9987954562051724
			 when "0011111001" => Y <= "000000011111101110011111001111100111111110"; -- Argumento 249( 1.5278448647340985 Radianes) Función 0.9990777277526454
			 when "0011111010" => Y <= "000000011111101110011111001111100111111001"; -- Argumento 250( 1.533980787885641 Radianes) Función 0.9993223845883495
			 when "0011111011" => Y <= "000000011111101110011111001111100111011011"; -- Argumento 251( 1.5401167110371838 Radianes) Función 0.9995294175010931
			 when "0011111100" => Y <= "000000011111101110011111001111100110011111"; -- Argumento 252( 1.5462526341887264 Radianes) Función 0.9996988186962042
			 when "0011111101" => Y <= "000000011111101110011111001111100111111111"; -- Argumento 253( 1.552388557340269 Radianes) Función 0.9998305817958234
			 when "0011111110" => Y <= "000000011111101110011111001111100111110011"; -- Argumento 254( 1.5585244804918115 Radianes) Función 0.9999247018391445
			 when "0011111111" => Y <= "000000011111101110011111001111100111110011"; -- Argumento 255( 1.564660403643354 Radianes) Función 0.9999811752826011
			 when "0100000000" => Y <= "000000001100001111110111111011111101111110"; -- Argumento 256( 1.5707963267948966 Radianes) Función 1.0
			 when "0100000001" => Y <= "000000011111101110011111001111100111110011"; -- Argumento 257( 1.576932249946439 Radianes) Función 0.9999811752826011
			 when "0100000010" => Y <= "000000011111101110011111001111100111110011"; -- Argumento 258( 1.5830681730979816 Radianes) Función 0.9999247018391445
			 when "0100000011" => Y <= "000000011111101110011111001111100111111111"; -- Argumento 259( 1.5892040962495242 Radianes) Función 0.9998305817958234
			 when "0100000100" => Y <= "000000011111101110011111001111100110011111"; -- Argumento 260( 1.5953400194010667 Radianes) Función 0.9996988186962042
			 when "0100000101" => Y <= "000000011111101110011111001111100111011011"; -- Argumento 261( 1.6014759425526093 Radianes) Función 0.9995294175010931
			 when "0100000110" => Y <= "000000011111101110011111001111100111111001"; -- Argumento 262( 1.607611865704152 Radianes) Función 0.9993223845883495
			 when "0100000111" => Y <= "000000011111101110011111001111100111111110"; -- Argumento 263( 1.6137477888556946 Radianes) Función 0.9990777277526454
			 when "0100001000" => Y <= "000000011111101110011111001111111111110001"; -- Argumento 264( 1.6198837120072371 Radianes) Función 0.9987954562051724
			 when "0100001001" => Y <= "000000011111101110011111001111111110110011"; -- Argumento 265( 1.6260196351587797 Radianes) Función 0.9984755805732948
			 when "0100001010" => Y <= "000000011111101110011111001111111110110000"; -- Argumento 266( 1.6321555583103222 Radianes) Función 0.9981181129001492
			 when "0100001011" => Y <= "000000011111101110011111001111100011110001"; -- Argumento 267( 1.6382914814618648 Radianes) Función 0.9977230666441916
			 when "0100001100" => Y <= "000000011111101110011111001111100011001101"; -- Argumento 268( 1.6444274046134073 Radianes) Función 0.9972904566786902
			 when "0100001101" => Y <= "000000011111101110011111001100111111111111"; -- Argumento 269( 1.6505633277649499 Radianes) Función 0.9968202992911657
			 when "0100001110" => Y <= "000000011111101110011111001100111111111001"; -- Argumento 270( 1.6566992509164924 Radianes) Función 0.996312612182778
			 when "0100001111" => Y <= "000000011111101110011111001110110111110001"; -- Argumento 271( 1.662835174068035 Radianes) Función 0.9957674144676598
			 when "0100010000" => Y <= "000000011111101110011111001110110110110000"; -- Argumento 272( 1.6689710972195777 Radianes) Función 0.9951847266721969
			 when "0100010001" => Y <= "000000011111101110011111001101100111011011"; -- Argumento 273( 1.6751070203711202 Radianes) Función 0.9945645707342554
			 when "0100010010" => Y <= "000000011111101110011111001111110011110011"; -- Argumento 274( 1.6812429435226628 Radianes) Función 0.9939069700023561
			 when "0100010011" => Y <= "000000011111101110011111001111110011001101"; -- Argumento 275( 1.6873788666742053 Radianes) Función 0.9932119492347945
			 when "0100010100" => Y <= "000000011111101110011111001110011010110011"; -- Argumento 276( 1.6935147898257479 Radianes) Función 0.99247953459871
			 when "0100010101" => Y <= "000000011111101110011111001101100001110001"; -- Argumento 277( 1.6996507129772904 Radianes) Función 0.9917097536690995
			 when "0100010110" => Y <= "000000011111101110011111001111111101110011"; -- Argumento 278( 1.705786636128833 Radianes) Función 0.99090263542778
			 when "0100010111" => Y <= "000000011111101110011111001111111101111110"; -- Argumento 279( 1.7119225592803755 Radianes) Función 0.9900582102622971
			 when "0100011000" => Y <= "000000011111101110011111111111100110110000"; -- Argumento 280( 1.718058482431918 Radianes) Función 0.989176509964781
			 when "0100011001" => Y <= "000000011111101110011111111111111111001101"; -- Argumento 281( 1.7241944055834606 Radianes) Función 0.9882575677307495
			 when "0100011010" => Y <= "000000011111101110011111111111100011111001"; -- Argumento 282( 1.7303303287350031 Radianes) Función 0.9873014181578584
			 when "0100011011" => Y <= "000000011111101110011111111100111111111001"; -- Argumento 283( 1.736466251886546 Radianes) Función 0.9863080972445987
			 when "0100011100" => Y <= "000000011111101110011111111110110111001101"; -- Argumento 284( 1.7426021750380885 Radianes) Función 0.9852776423889412
			 when "0100011101" => Y <= "000000011111101110011111111101100111001101"; -- Argumento 285( 1.748738098189631 Radianes) Función 0.984210092386929
			 when "0100011110" => Y <= "000000011111101110011111111111110010110000"; -- Argumento 286( 1.7548740213411735 Radianes) Función 0.9831054874312163
			 when "0100011111" => Y <= "000000011111101110011111111101100001110011"; -- Argumento 287( 1.761009944492716 Radianes) Función 0.9819638691095552
			 when "0100100000" => Y <= "000000011111101110011111111111111101110001"; -- Argumento 288( 1.7671458676442586 Radianes) Función 0.9807852804032304
			 when "0100100001" => Y <= "000000011111101110011111000111100111011011"; -- Argumento 289( 1.7732817907958012 Radianes) Función 0.9795697656854405
			 when "0100100010" => Y <= "000000011111101110011111000111111111111001"; -- Argumento 290( 1.7794177139473437 Radianes) Función 0.9783173707196277
			 when "0100100011" => Y <= "000000011111101110011111000111100011111110"; -- Argumento 291( 1.7855536370988863 Radianes) Función 0.9770281426577544
			 when "0100100100" => Y <= "000000011111101110011111000110110111110001"; -- Argumento 292( 1.7916895602504288 Radianes) Función 0.9757021300385286
			 when "0100100101" => Y <= "000000011111101110011111000101100111111001"; -- Argumento 293( 1.7978254834019713 Radianes) Función 0.9743393827855759
			 when "0100100110" => Y <= "000000011111101110011111000110011011110011"; -- Argumento 294( 1.8039614065535141 Radianes) Función 0.9729399522055602
			 when "0100100111" => Y <= "000000011111101110011111000101100001011011"; -- Argumento 295( 1.8100973297050567 Radianes) Función 0.9715038909862518
			 when "0100101000" => Y <= "000000011111101110011111000111111101111110"; -- Argumento 296( 1.8162332528565992 Radianes) Función 0.970031253194544
			 when "0100101001" => Y <= "000000011111101110011001111111111111011011"; -- Argumento 297( 1.8223691760081417 Radianes) Función 0.9685220942744174
			 when "0100101010" => Y <= "000000011111101110011001111100111111110011"; -- Argumento 298( 1.8285050991596843 Radianes) Función 0.9669764710448521
			 when "0100101011" => Y <= "000000011111101110011001111110110111111001"; -- Argumento 299( 1.8346410223112268 Radianes) Función 0.9653944416976894
			 when "0100101100" => Y <= "000000011111101110011001111111110011110001"; -- Argumento 300( 1.8407769454627694 Radianes) Función 0.9637760657954398
			 when "0100101101" => Y <= "000000011111101110011001111110011010110000"; -- Argumento 301( 1.846912868614312 Radianes) Función 0.9621214042690416
			 when "0100101110" => Y <= "000000011111101110011001111111111100110011"; -- Argumento 302( 1.8530487917658545 Radianes) Función 0.9604305194155659
			 when "0100101111" => Y <= "000000011111101110011101101111111111110001"; -- Argumento 303( 1.859184714917397 Radianes) Función 0.9587034748958716
			 when "0100110000" => Y <= "000000011111101110011101101100111111110011"; -- Argumento 304( 1.8653206380689396 Radianes) Función 0.9569403357322089
			 when "0100110001" => Y <= "000000011111101110011101101110110110110000"; -- Argumento 305( 1.8714565612204823 Radianes) Función 0.9551411683057707
			 when "0100110010" => Y <= "000000011111101110011101101111110011111001"; -- Argumento 306( 1.8775924843720249 Radianes) Función 0.9533060403541939
			 when "0100110011" => Y <= "000000011111101110011101101101100000110011"; -- Argumento 307( 1.8837284075235674 Radianes) Función 0.9514350209690083
			 when "0100110100" => Y <= "000000011111101110011011001111100111011011"; -- Argumento 308( 1.88986433067511 Radianes) Función 0.9495281805930367
			 when "0100110101" => Y <= "000000011111101110011011001111100011011011"; -- Argumento 309( 1.8960002538266525 Radianes) Función 0.9475855910177412
			 when "0100110110" => Y <= "000000011111101110011011001110110110011111"; -- Argumento 310( 1.902136176978195 Radianes) Función 0.9456073253805214
			 when "0100110111" => Y <= "000000011111101110011011001111110011011011"; -- Argumento 311( 1.9082721001297376 Radianes) Función 0.9435934581619604
			 when "0100111000" => Y <= "000000011111101110011011001101100001011011"; -- Argumento 312( 1.9144080232812801 Radianes) Función 0.9415440651830208
			 when "0100111001" => Y <= "000000011111101110011111100111100110110011"; -- Argumento 313( 1.9205439464328227 Radianes) Función 0.9394592236021899
			 when "0100111010" => Y <= "000000011111101110011111100111100011111001"; -- Argumento 314( 1.9266798695843652 Radianes) Función 0.937339011912575
			 when "0100111011" => Y <= "000000011111101110011111100110110110110000"; -- Argumento 315( 1.932815792735908 Radianes) Función 0.9351835099389476
			 when "0100111100" => Y <= "000000011111101110011111100110011011110011"; -- Argumento 316( 1.9389517158874505 Radianes) Función 0.9329927988347388
			 when "0100111101" => Y <= "000000011111101110011111100111111101110001"; -- Argumento 317( 1.945087639038993 Radianes) Función 0.9307669610789837
			 when "0100111110" => Y <= "000000011111101110011100110111111111011011"; -- Argumento 318( 1.9512235621905356 Radianes) Función 0.9285060804732156
			 when "0100111111" => Y <= "000000011111101110011100110100111111001101"; -- Argumento 319( 1.9573594853420782 Radianes) Función 0.9262102421383114
			 when "0101000000" => Y <= "000000011111101110011100110111110011111111"; -- Argumento 320( 1.9634954084936207 Radianes) Función 0.9238795325112867
			 when "0101000001" => Y <= "000000011111101110011100110101100001011011"; -- Argumento 321( 1.9696313316451632 Radianes) Función 0.921514039342042
			 when "0101000010" => Y <= "000000011111101110011011000011100110110000"; -- Argumento 322( 1.9757672547967058 Radianes) Función 0.9191138516900578
			 when "0101000011" => Y <= "000000011111101110011011000000111110011111"; -- Argumento 323( 1.9819031779482483 Radianes) Función 0.9166790599210427
			 when "0101000100" => Y <= "000000011111101110011011000001100111001101"; -- Argumento 324( 1.9880391010997909 Radianes) Función 0.9142097557035307
			 when "0101000101" => Y <= "000000011111101110011011000001100001110001"; -- Argumento 325( 1.9941750242513334 Radianes) Función 0.9117060320054299
			 when "0101000110" => Y <= "000000011111101110011111111011100110110000"; -- Argumento 326( 2.000310947402876 Radianes) Función 0.9091679830905225
			 when "0101000111" => Y <= "000000011111101110011111111000111111011011"; -- Argumento 327( 2.0064468705544187 Radianes) Función 0.9065957045149153
			 when "0101001000" => Y <= "000000011111101110011111111011110011110011"; -- Argumento 328( 2.012582793705961 Radianes) Función 0.9039892931234434
			 when "0101001001" => Y <= "000000011111101110011111111001100001111001"; -- Argumento 329( 2.018718716857504 Radianes) Función 0.901348847046022
			 when "0101001010" => Y <= "000000011111101111111111001111111110011111"; -- Argumento 330( 2.024854640009046 Radianes) Función 0.8986744656939539
			 when "0101001011" => Y <= "000000011111101111111111001110110111110011"; -- Argumento 331( 2.030990563160589 Radianes) Función 0.8959662497561852
			 when "0101001100" => Y <= "000000011111101111111111001111110011001101"; -- Argumento 332( 2.0371264863121317 Radianes) Función 0.8932243011955152
			 when "0101001101" => Y <= "000000011111101111111111001111111100110011"; -- Argumento 333( 2.043262409463674 Radianes) Función 0.890448723244758
			 when "0101001110" => Y <= "000000011111101111111111111111100010011111"; -- Argumento 334( 2.0493983326152168 Radianes) Función 0.8876396204028539
			 when "0101001111" => Y <= "000000011111101111111111111101100111110001"; -- Argumento 335( 2.055534255766759 Radianes) Función 0.8847970984309379
			 when "0101010000" => Y <= "000000011111101111111111111101100001110011"; -- Argumento 336( 2.061670178918302 Radianes) Función 0.881921264348355
			 when "0101010001" => Y <= "000000011111101111111111000111100111111110"; -- Argumento 337( 2.067806102069844 Radianes) Función 0.8790122264286335
			 when "0101010010" => Y <= "000000011111101111111111000100111111111110"; -- Argumento 338( 2.073942025221387 Radianes) Función 0.8760700941954066
			 when "0101010011" => Y <= "000000011111101111111111000111110011111110"; -- Argumento 339( 2.0800779483729293 Radianes) Función 0.8730949784182902
			 when "0101010100" => Y <= "000000011111101111111111000111111101111110"; -- Argumento 340( 2.086213871524472 Radianes) Función 0.8700869911087115
			 when "0101010101" => Y <= "000000011111101111111001111111100011111110"; -- Argumento 341( 2.0923497946760143 Radianes) Función 0.8670462455156928
			 when "0101010110" => Y <= "000000011111101111111001111111110011110011"; -- Argumento 342( 2.098485717827557 Radianes) Función 0.8639728561215868
			 when "0101010111" => Y <= "000000011111101111111001111111111101111111"; -- Argumento 343( 2.1046216409791 Radianes) Función 0.8608669386377672
			 when "0101011000" => Y <= "000000011111101111111101101111100011110001"; -- Argumento 344( 2.110757564130642 Radianes) Función 0.8577286100002721
			 when "0101011001" => Y <= "000000011111101111111101101101100111011011"; -- Argumento 345( 2.116893487282185 Radianes) Función 0.8545579883654005
			 when "0101011010" => Y <= "000000011111101111111101101101100001111001"; -- Argumento 346( 2.1230294104337273 Radianes) Función 0.8513551931052653
			 when "0101011011" => Y <= "000000011111101111111011001111111110110000"; -- Argumento 347( 2.12916533358527 Radianes) Función 0.8481203448032972
			 when "0101011100" => Y <= "000000011111101111111011001101100111111111"; -- Argumento 348( 2.1353012567368124 Radianes) Función 0.8448535652497072
			 when "0101011101" => Y <= "000000011111101111111011001101100001011011"; -- Argumento 349( 2.141437179888355 Radianes) Función 0.8415549774368984
			 when "0101011110" => Y <= "000000011111101111111111100111111111001101"; -- Argumento 350( 2.1475731030398975 Radianes) Función 0.8382247055548382
			 when "0101011111" => Y <= "000000011111101111111111100101100111111111"; -- Argumento 351( 2.1537090261914402 Radianes) Función 0.8348628749863801
			 when "0101100000" => Y <= "000000011111101111111111100101100000110011"; -- Argumento 352( 2.1598449493429825 Radianes) Función 0.8314696123025455
			 when "0101100001" => Y <= "000000011111101111111100110111111111111110"; -- Argumento 353( 2.1659808724945253 Radianes) Función 0.8280450452577558
			 when "0101100010" => Y <= "000000011111101111111100110101100111011011"; -- Argumento 354( 2.172116795646068 Radianes) Función 0.8245893027850253
			 when "0101100011" => Y <= "000000011111101111111100110101100000110000"; -- Argumento 355( 2.1782527187976104 Radianes) Función 0.8211025149911048
			 when "0101100100" => Y <= "000000011111101111111011000011100011011011"; -- Argumento 356( 2.184388641949153 Radianes) Función 0.8175848131515837
			 when "0101100101" => Y <= "000000011111101111111011000001100111111110"; -- Argumento 357( 2.1905245651006955 Radianes) Función 0.8140363297059485
			 when "0101100110" => Y <= "000000011111101111111011000011111100110011"; -- Argumento 358( 2.1966604882522383 Radianes) Función 0.8104571982525948
			 when "0101100111" => Y <= "000000011111101111111111111000111111111111"; -- Argumento 359( 2.2027964114037806 Radianes) Función 0.8068475535437994
			 when "0101101000" => Y <= "000000011111101111111111111011110011001101"; -- Argumento 360( 2.2089323345553233 Radianes) Función 0.8032075314806449
			 when "0101101001" => Y <= "000000011111101110001111001111100111011011"; -- Argumento 361( 2.2150682577068657 Radianes) Función 0.7995372691079052
			 when "0101101010" => Y <= "000000011111101110001111001110110111111111"; -- Argumento 362( 2.2212041808584084 Radianes) Función 0.7958369046088836
			 when "0101101011" => Y <= "000000011111101110001111001110011010110000"; -- Argumento 363( 2.227340104009951 Radianes) Función 0.7921065773002123
			 when "0101101100" => Y <= "000000011111101110001111111111111111111001"; -- Argumento 364( 2.2334760271614935 Radianes) Función 0.7883464276266063
			 when "0101101101" => Y <= "000000011111101110001111111101100111011011"; -- Argumento 365( 2.2396119503130363 Radianes) Función 0.7845565971555752
			 when "0101101110" => Y <= "000000011111101110001111111111111101110001"; -- Argumento 366( 2.2457478734645786 Radianes) Función 0.7807372285720946
			 when "0101101111" => Y <= "000000011111101110001111000100111111111111"; -- Argumento 367( 2.2518837966161214 Radianes) Función 0.7768884656732324
			 when "0101110000" => Y <= "000000011111101110001111000111110011111110"; -- Argumento 368( 2.2580197197676637 Radianes) Función 0.7730104533627371
			 when "0101110001" => Y <= "000000011111101110001001111111100110110000"; -- Argumento 369( 2.2641556429192065 Radianes) Función 0.7691033376455797
			 when "0101110010" => Y <= "000000011111101110001001111110110110110000"; -- Argumento 370( 2.270291566070749 Radianes) Función 0.7651672656224591
			 when "0101110011" => Y <= "000000011111101110001001111101100001001101"; -- Argumento 371( 2.2764274892222915 Radianes) Función 0.7612023854842619
			 when "0101110100" => Y <= "000000011111101110001101101111100011001101"; -- Argumento 372( 2.282563412373834 Radianes) Función 0.7572088465064848
			 when "0101110101" => Y <= "000000011111101110001101101111110010110000"; -- Argumento 373( 2.2886993355253766 Radianes) Función 0.7531867990436125
			 when "0101110110" => Y <= "000000011111101110001011001111100110110000"; -- Argumento 374( 2.2948352586769194 Radianes) Función 0.7491363945234593
			 when "0101110111" => Y <= "000000011111101110001011001110110111111110"; -- Argumento 375( 2.3009711818284617 Radianes) Función 0.7450577854414661
			 when "0101111000" => Y <= "000000011111101110001011001111111101110011"; -- Argumento 376( 2.3071071049800045 Radianes) Función 0.7409511253549591
			 when "0101111001" => Y <= "000000011111101110001111100100111111111111"; -- Argumento 377( 2.313243028131547 Radianes) Función 0.73681656887737
			 when "0101111010" => Y <= "000000011111101110001111100110011010011111"; -- Argumento 378( 2.3193789512830896 Radianes) Función 0.7326542716724128
			 when "0101111011" => Y <= "000000011111101110001100110111111110110011"; -- Argumento 379( 2.325514874434632 Radianes) Función 0.7284643904482253
			 when "0101111100" => Y <= "000000011111101110001100110101100111001101"; -- Argumento 380( 2.3316507975861747 Radianes) Función 0.724247082951467
			 when "0101111101" => Y <= "000000011111101110001100110111111101111110"; -- Argumento 381( 2.337786720737717 Radianes) Función 0.7200025079613818
			 when "0101111110" => Y <= "000000011111101110001011000010110111110001"; -- Argumento 382( 2.3439226438892597 Radianes) Función 0.7157308252838187
			 when "0101111111" => Y <= "000000011111101110001011000001100000110011"; -- Argumento 383( 2.350058567040802 Radianes) Función 0.7114321957452167
			 when "0110000000" => Y <= "000000011111101110001111111011100010110000"; -- Argumento 384( 2.356194490192345 Radianes) Función 0.7071067811865476
			 when "0110000001" => Y <= "000000011111101110001111111010011011110001"; -- Argumento 385( 2.3623304133438876 Radianes) Función 0.7027547444572252
			 when "0110000010" => Y <= "000000011111100011111111001111111111111001"; -- Argumento 386( 2.36846633649543 Radianes) Función 0.6983762494089729
			 when "0110000011" => Y <= "000000011111100011111111001111110011110011"; -- Argumento 387( 2.3746022596469727 Radianes) Función 0.693971460889654
			 when "0110000100" => Y <= "000000011111100011111111111111100111011011"; -- Argumento 388( 2.380738182798515 Radianes) Función 0.689540544737067
			 when "0110000101" => Y <= "000000011111100011111111111110110111111110"; -- Argumento 389( 2.386874105950058 Radianes) Función 0.6850836677727004
			 when "0110000110" => Y <= "000000011111100011111111111111111100011111"; -- Argumento 390( 2.3930100291016 Radianes) Función 0.6806009977954532
			 when "0110000111" => Y <= "000000011111100011111111000100111111111110"; -- Argumento 391( 2.399145952253143 Radianes) Función 0.6760927035753159
			 when "0110001000" => Y <= "000000011111100011111111000101100001011011"; -- Argumento 392( 2.405281875404685 Radianes) Función 0.6715589548470186
			 when "0110001001" => Y <= "000000011111100011111001111100111111110011"; -- Argumento 393( 2.411417798556228 Radianes) Función 0.6669999223036376
			 when "0110001010" => Y <= "000000011111100011111001111110011010110011"; -- Argumento 394( 2.4175537217077703 Radianes) Función 0.662415777590172
			 when "0110001011" => Y <= "000000011111100011111101101111100011111111"; -- Argumento 395( 2.423689644859313 Radianes) Función 0.6578066932970787
			 when "0110001100" => Y <= "000000011111100011111101101111110010110000"; -- Argumento 396( 2.429825568010856 Radianes) Función 0.6531728429537766
			 when "0110001101" => Y <= "000000011111100011111011001111111111011011"; -- Argumento 397( 2.435961491162398 Radianes) Función 0.6485144010221126
			 when "0110001110" => Y <= "000000011111100011111011001111110011111111"; -- Argumento 398( 2.442097414313941 Radianes) Función 0.6438315428897914
			 when "0110001111" => Y <= "000000011111100011111111100111100110110000"; -- Argumento 399( 2.448233337465483 Radianes) Función 0.6391244448637758
			 when "0110010000" => Y <= "000000011111100011111111100101100111111001"; -- Argumento 400( 2.454369260617026 Radianes) Función 0.6343932841636455
			 when "0110010001" => Y <= "000000011111100011111100110111100110011111"; -- Argumento 401( 2.4605051837685683 Radianes) Función 0.6296382389149272
			 when "0110010010" => Y <= "000000011111100011111100110101100111111111"; -- Argumento 402( 2.466641106920111 Radianes) Función 0.6248594881423863
			 when "0110010011" => Y <= "000000011111100011111100110111111101111110"; -- Argumento 403( 2.4727770300716534 Radianes) Función 0.6200572117632894
			 when "0110010100" => Y <= "000000011111100011111011000010110111001101"; -- Argumento 404( 2.478912953223196 Radianes) Función 0.6152315905806269
			 when "0110010101" => Y <= "000000011111100011111011000011111101111001"; -- Argumento 405( 2.4850488763747385 Radianes) Función 0.6103828062763097
			 when "0110010110" => Y <= "000000011111100011111111111010110111011011"; -- Argumento 406( 2.4911847995262812 Radianes) Función 0.6055110414043255
			 when "0110010111" => Y <= "000000011111100011111111111011111100011111"; -- Argumento 407( 2.497320722677824 Radianes) Función 0.6006164793838689
			 when "0110011000" => Y <= "000000011111101011011111001110110110011111"; -- Argumento 408( 2.5034566458293663 Radianes) Función 0.5956993044924335
			 when "0110011001" => Y <= "000000011111101011011111001111111101110001"; -- Argumento 409( 2.509592568980909 Radianes) Función 0.5907597018588742
			 when "0110011010" => Y <= "000000011111101011011111111110110111110001"; -- Argumento 410( 2.5157284921324514 Radianes) Función 0.585797857456439
			 when "0110011011" => Y <= "000000011111101011011111111111111101111111"; -- Argumento 411( 2.521864415283994 Radianes) Función 0.5808139580957645
			 when "0110011100" => Y <= "000000011111101011011111000110110111111111"; -- Argumento 412( 2.5280003384355365 Radianes) Función 0.5758081914178454
			 when "0110011101" => Y <= "000000011111101011011111000111111101110001"; -- Argumento 413( 2.5341362615870793 Radianes) Función 0.5707807458869673
			 when "0110011110" => Y <= "000000011111101011011001111110110111110001"; -- Argumento 414( 2.5402721847386216 Radianes) Función 0.5657318107836135
			 when "0110011111" => Y <= "000000011111101011011001111111111100011111"; -- Argumento 415( 2.5464081078901644 Radianes) Función 0.560661576197336
			 when "0110100000" => Y <= "000000011111101011011101101110110111011011"; -- Argumento 416( 2.552544031041707 Radianes) Función 0.5555702330196021
			 when "0110100001" => Y <= "000000011111101011011101101111111100110011"; -- Argumento 417( 2.5586799541932495 Radianes) Función 0.5504579729366049
			 when "0110100010" => Y <= "000000011111101011011011001110110111111001"; -- Argumento 418( 2.564815877344792 Radianes) Función 0.5453249884220464
			 when "0110100011" => Y <= "000000011111101011011011001111111100110000"; -- Argumento 419( 2.5709518004963345 Radianes) Función 0.540171472729893
			 when "0110100100" => Y <= "000000011111101011011111100101100111110011"; -- Argumento 420( 2.5770877236478773 Radianes) Función 0.5349976198870972
			 when "0110100101" => Y <= "000000011111101011011100110111100111111111"; -- Argumento 421( 2.5832236467994196 Radianes) Función 0.5298036246862948
			 when "0110100110" => Y <= "000000011111101011011100110101100111011011"; -- Argumento 422( 2.5893595699509624 Radianes) Función 0.524589682678469
			 when "0110100111" => Y <= "000000011111101011011011000011100111111001"; -- Argumento 423( 2.5954954931025047 Radianes) Función 0.5193559901655898
			 when "0110101000" => Y <= "000000011111101011011011000001100110110000"; -- Argumento 424( 2.6016314162540475 Radianes) Función 0.5141027441932218
			 when "0110101001" => Y <= "000000011111101011011111111011111111111111"; -- Argumento 425( 2.60776733940559 Radianes) Función 0.5088301425431073
			 when "0110101010" => Y <= "000000011111101011011111111011110011011011"; -- Argumento 426( 2.6139032625571326 Radianes) Función 0.5035383837257176
			 when "0110101011" => Y <= "000000011111100110011111001111111111001101"; -- Argumento 427( 2.6200391857086753 Radianes) Función 0.49822766697278176
			 when "0110101100" => Y <= "000000011111100110011111001110011011111111"; -- Argumento 428( 2.6261751088602177 Radianes) Función 0.49289819222978415
			 when "0110101101" => Y <= "000000011111100110011111111111100011011011"; -- Argumento 429( 2.6323110320117604 Radianes) Función 0.4875501601484359
			 when "0110101110" => Y <= "000000011111100110011111111110011010110000"; -- Argumento 430( 2.6384469551633027 Radianes) Función 0.4821837720791229
			 when "0110101111" => Y <= "000000011111100110011111000100111111110001"; -- Argumento 431( 2.6445828783148455 Radianes) Función 0.4767992300633221
			 when "0110110000" => Y <= "000000011111100110011111000101100001111001"; -- Argumento 432( 2.650718801466388 Radianes) Función 0.4713967368259978
			 when "0110110001" => Y <= "000000011111100110011001111110110111110011"; -- Argumento 433( 2.6568547246179306 Radianes) Función 0.4659764957679662
			 when "0110110010" => Y <= "000000011111100110011001111111111101011011"; -- Argumento 434( 2.662990647769473 Radianes) Función 0.4605387109582402
			 when "0110110011" => Y <= "000000011111100110011101101110110111111110"; -- Argumento 435( 2.6691265709210157 Radianes) Función 0.4550835871263439
			 when "0110110100" => Y <= "000000011111100110011011001111100110011111"; -- Argumento 436( 2.675262494072558 Radianes) Función 0.4496113296546069
			 when "0110110101" => Y <= "000000011111100110011011001101100110110000"; -- Argumento 437( 2.6813984172241008 Radianes) Función 0.4441221445704293
			 when "0110110110" => Y <= "000000011111100110011111100111111110011111"; -- Argumento 438( 2.6875343403756435 Radianes) Función 0.43861623853852755
			 when "0110110111" => Y <= "000000011111100110011111100111110011111110"; -- Argumento 439( 2.693670263527186 Radianes) Función 0.43309381885315207
			 when "0110111000" => Y <= "000000011111100110011100110111100011011011"; -- Argumento 440( 2.6998061866787286 Radianes) Función 0.42755509343028203
			 when "0110111001" => Y <= "000000011111100110011100110110011011111110"; -- Argumento 441( 2.705942109830271 Radianes) Función 0.42200027079979985
			 when "0110111010" => Y <= "000000011111100110011011000000111110110011"; -- Argumento 442( 2.7120780329818137 Radianes) Función 0.41642956009763715
			 when "0110111011" => Y <= "000000011111100110011011000011111101111111"; -- Argumento 443( 2.718213956133356 Radianes) Función 0.41084317105790413
			 when "0110111100" => Y <= "000000011111100110011111111010110111001101"; -- Argumento 444( 2.724349879284899 Radianes) Función 0.40524131400498986
			 when "0110111101" => Y <= "000000011111101111001111001111100110011111"; -- Argumento 445( 2.730485802436441 Radianes) Función 0.39962419984564707
			 when "0110111110" => Y <= "000000011111101111001111001111110011110011"; -- Argumento 446( 2.736621725587984 Radianes) Función 0.39399204006104815
			 when "0110111111" => Y <= "000000011111101111001111111111111111111001"; -- Argumento 447( 2.742757648739526 Radianes) Función 0.3883450466988266
			 when "0111000000" => Y <= "000000011111101111001111111110011010011111"; -- Argumento 448( 2.748893571891069 Radianes) Función 0.38268343236508984
			 when "0111000001" => Y <= "000000011111101111001111000111100011111110"; -- Argumento 449( 2.7550294950426117 Radianes) Función 0.37700741021641815
			 when "0111000010" => Y <= "000000011111101111001111000101100001111001"; -- Argumento 450( 2.761165418194154 Radianes) Función 0.37131719395183765
			 when "0111000011" => Y <= "000000011111101111001001111110110110011111"; -- Argumento 451( 2.767301341345697 Radianes) Función 0.3656129978047738
			 when "0111000100" => Y <= "000000011111101111001101101111100111111111"; -- Argumento 452( 2.773437264497239 Radianes) Función 0.35989503653498833
			 when "0111000101" => Y <= "000000011111101111001101101101100110110000"; -- Argumento 453( 2.779573187648782 Radianes) Función 0.35416352542049034
			 when "0111000110" => Y <= "000000011111101111001011001111111110110011"; -- Argumento 454( 2.7857091108003242 Radianes) Función 0.3484186802494348
			 when "0111000111" => Y <= "000000011111101111001011001110011010011111"; -- Argumento 455( 2.791845033951867 Radianes) Función 0.34266071731199443
			 when "0111001000" => Y <= "000000011111101111001111100100111111111111"; -- Argumento 456( 2.7979809571034093 Radianes) Función 0.3368898533922203
			 when "0111001001" => Y <= "000000011111101111001111100101100000110000"; -- Argumento 457( 2.804116880254952 Radianes) Función 0.3311063057598765
			 when "0111001010" => Y <= "000000011111101111001100110110110111111001"; -- Argumento 458( 2.8102528034064944 Radianes) Función 0.3253102921622632
			 when "0111001011" => Y <= "000000011111101111001011000011100111011011"; -- Argumento 459( 2.816388726558037 Radianes) Función 0.3195020308160158
			 when "0111001100" => Y <= "000000011111101111001011000011110010011111"; -- Argumento 460( 2.82252464970958 Radianes) Función 0.3136817403988914
			 when "0111001101" => Y <= "000000011111101111001111111011100011111111"; -- Argumento 461( 2.8286605728611223 Radianes) Función 0.30784964004153503
			 when "0111001110" => Y <= "000000011111101111001111111010011011111110"; -- Argumento 462( 2.834796496012665 Radianes) Función 0.30200594931922803
			 when "0111001111" => Y <= "000000011111101001101111001100111110110000"; -- Argumento 463( 2.8409324191642074 Radianes) Función 0.296150888243624
			 when "0111010000" => Y <= "000000011111101001101111001111111101001101"; -- Argumento 464( 2.84706834231575 Radianes) Función 0.29028467725446233
			 when "0111010001" => Y <= "000000011111101001101111111101100110110011"; -- Argumento 465( 2.8532042654672924 Radianes) Función 0.28440753721127204
			 when "0111010010" => Y <= "000000011111101001101111000111111111011011"; -- Argumento 466( 2.859340188618835 Radianes) Función 0.2785196893850531
			 when "0111010011" => Y <= "000000011111101001101111000110011010011111"; -- Argumento 467( 2.8654761117703775 Radianes) Función 0.27262135544994925
			 when "0111010100" => Y <= "000000011111101001101001111100111111110001"; -- Argumento 468( 2.8716120349219203 Radianes) Función 0.2667127574748985
			 when "0111010101" => Y <= "000000011111101001101001111111111101110001"; -- Argumento 469( 2.8777479580734626 Radianes) Función 0.26079411791527585
			 when "0111010110" => Y <= "000000011111101001101101101101100111111111"; -- Argumento 470( 2.8838838812250054 Radianes) Función 0.2548656596045147
			 when "0111010111" => Y <= "000000011111101001101011001111111111110011"; -- Argumento 471( 2.890019804376548 Radianes) Función 0.2489276057457201
			 when "0111011000" => Y <= "000000011111101001101011001110011011110011"; -- Argumento 472( 2.8961557275280905 Radianes) Función 0.24298017990326404
			 when "0111011001" => Y <= "000000011111101001101111100111100011111110"; -- Argumento 473( 2.9022916506796332 Radianes) Función 0.23702360599436717
			 when "0111011010" => Y <= "000000011111101001101111100101100001111110"; -- Argumento 474( 2.9084275738311756 Radianes) Función 0.2310581082806713
			 when "0111011011" => Y <= "000000011111101001101100110110110111111110"; -- Argumento 475( 2.9145634969827183 Radianes) Función 0.22508391135979283
			 when "0111011100" => Y <= "000000011111101001101011000011100110110000"; -- Argumento 476( 2.9206994201342606 Radianes) Función 0.21910124015687002
			 when "0111011101" => Y <= "000000011111101001101011000011110010110000"; -- Argumento 477( 2.9268353432858034 Radianes) Función 0.21311031991609142
			 when "0111011110" => Y <= "000000011111101001101111111011100010110000"; -- Argumento 478( 2.9329712664373457 Radianes) Función 0.20711137619221884
			 when "0111011111" => Y <= "000000011111101001101111111001100000110000"; -- Argumento 479( 2.9391071895888885 Radianes) Función 0.20110463484209198
			 when "0111100000" => Y <= "000000011111100110000111001110110111111110"; -- Argumento 480( 2.945243112740431 Radianes) Función 0.19509032201612858
			 when "0111100001" => Y <= "000000011111100110000111111111100111111110"; -- Argumento 481( 2.9513790358919736 Radianes) Función 0.18906866414980633
			 when "0111100010" => Y <= "000000011111100110000111111111110011111110"; -- Argumento 482( 2.9575149590435164 Radianes) Función 0.1830398879551409
			 when "0111100011" => Y <= "000000011111100110000111000111100011111110"; -- Argumento 483( 2.9636508821950587 Radianes) Función 0.17700422041214892
			 when "0111100100" => Y <= "000000011111100110000111000111111101110011"; -- Argumento 484( 2.9697868053466014 Radianes) Función 0.1709618887603012
			 when "0111100101" => Y <= "000000011111100110000001111101100111110011"; -- Argumento 485( 2.9759227284981438 Radianes) Función 0.16491312048997012
			 when "0111100110" => Y <= "000000011111100110000101101111111111111111"; -- Argumento 486( 2.9820586516496865 Radianes) Función 0.15885814333386145
			 when "0111100111" => Y <= "000000011111100110000101101110011011110001"; -- Argumento 487( 2.988194574801229 Radianes) Función 0.15279718525844369
			 when "0111101000" => Y <= "000000011111100110000011001100111111110001"; -- Argumento 488( 2.9943304979527716 Radianes) Función 0.1467304744553618
			 when "0111101001" => Y <= "000000011111100110000011001111111100011111"; -- Argumento 489( 3.000466421104314 Radianes) Función 0.14065823933284952
			 when "0111101010" => Y <= "000000011111100110000111100101100111011011"; -- Argumento 490( 3.0066023442558567 Radianes) Función 0.13458070850712628
			 when "0111101011" => Y <= "000000011111100110000100110111111110110011"; -- Argumento 491( 3.0127382674073995 Radianes) Función 0.12849811079379306
			 when "0111101100" => Y <= "000000011111100110000100110110011010110011"; -- Argumento 492( 3.018874190558942 Radianes) Función 0.12241067519921635
			 when "0111101101" => Y <= "000000011111100110000011000000111111111001"; -- Argumento 493( 3.0250101137104846 Radianes) Función 0.11631863091190471
			 when "0111101110" => Y <= "000000011111100110000011000011111101001101"; -- Argumento 494( 3.031146036862027 Radianes) Función 0.11022220729388325
			 when "0111101111" => Y <= "000000011111100110000111111001100110110000"; -- Argumento 495( 3.0372819600135696 Radianes) Función 0.10412163387205457
			 when "0111110000" => Y <= "000000011111101111110111001111111111111110"; -- Argumento 496( 3.043417883165112 Radianes) Función 0.09801714032956084
			 when "0111110001" => Y <= "000000011111101111110111001101100001110011"; -- Argumento 497( 3.0495538063166547 Radianes) Función 0.09190895649713277
			 when "0111110010" => Y <= "000000011111101111110111111110110111110001"; -- Argumento 498( 3.055689729468197 Radianes) Función 0.08579731234444016
			 when "0111110011" => Y <= "000000011111101111110111000111100110011111"; -- Argumento 499( 3.06182565261974 Radianes) Función 0.0796824379714302
			 when "0111110100" => Y <= "000000011111101111110111000111110011011011"; -- Argumento 500( 3.067961575771282 Radianes) Función 0.07356456359966775
			 when "0111110101" => Y <= "000000011111101111110001111111100010110011"; -- Argumento 501( 3.074097498922825 Radianes) Función 0.06744391956366418
			 when "0111110110" => Y <= "000000011111101111110001111101100001111001"; -- Argumento 502( 3.0802334220743677 Radianes) Función 0.061320736302208495
			 when "0111110111" => Y <= "000000011111101111110101101110110110110000"; -- Argumento 503( 3.08636934522591 Radianes) Función 0.055195244349690094
			 when "0111111000" => Y <= "000000011111101111110011001111100111111110"; -- Argumento 504( 3.0925052683774528 Radianes) Función 0.04906767432741797
			 when "0111111001" => Y <= "000000011111101111110011001110011011110011"; -- Argumento 505( 3.098641191528995 Radianes) Función 0.04293825693494102
			 when "0111111010" => Y <= "000000011111101111110111100100111111111111"; -- Argumento 506( 3.104777114680538 Radianes) Función 0.03680722294135883
			 when "0111111011" => Y <= "000000011111101111110111100111111100011111"; -- Argumento 507( 3.11091303783208 Radianes) Función 0.030674803176636865
			 when "0111111100" => Y <= "000000011111101111110100110101100111011011"; -- Argumento 508( 3.117048960983623 Radianes) Función 0.024541228522912326
			 when "0111111101" => Y <= "000000011111101111110011000011111110110011"; -- Argumento 509( 3.1231848841351653 Radianes) Función 0.0184067299058051
			 when "0111111110" => Y <= "000000011111101111110011000010011011001101"; -- Argumento 510( 3.129320807286708 Radianes) Función 0.012271538285720007
			 when "0111111111" => Y <= "000000011111101111110111111000111110110000"; -- Argumento 511( 3.1354567304382504 Radianes) Función 0.006135884649154799
			 when "1000000000" => Y <= "000000011111101111110111111011111101111110"; -- Argumento 512( 3.141592653589793 Radianes) Función 1.2246467991473532e-16
			 when "1000000001" => Y <= "000000111111101111110111111000111110110000"; -- Argumento 513( 3.147728576741336 Radianes) Función -0.006135884649154554
			 when "1000000010" => Y <= "000000111111101111110011000010011011001101"; -- Argumento 514( 3.153864499892878 Radianes) Función -0.01227153828571976
			 when "1000000011" => Y <= "000000111111101111110011000011111110110011"; -- Argumento 515( 3.160000423044421 Radianes) Función -0.01840672990580486
			 when "1000000100" => Y <= "000000111111101111110100110101100111011011"; -- Argumento 516( 3.1661363461959633 Radianes) Función -0.024541228522912083
			 when "1000000101" => Y <= "000000111111101111110111100111111100011111"; -- Argumento 517( 3.172272269347506 Radianes) Función -0.030674803176636622
			 when "1000000110" => Y <= "000000111111101111110111100100111111111111"; -- Argumento 518( 3.1784081924990484 Radianes) Función -0.03680722294135858
			 when "1000000111" => Y <= "000000111111101111110011001110011011110011"; -- Argumento 519( 3.184544115650591 Radianes) Función -0.04293825693494077
			 when "1000001000" => Y <= "000000111111101111110011001111100111111110"; -- Argumento 520( 3.1906800388021335 Radianes) Función -0.049067674327417724
			 when "1000001001" => Y <= "000000111111101111110101101110110110110000"; -- Argumento 521( 3.1968159619536762 Radianes) Función -0.05519524434968985
			 when "1000001010" => Y <= "000000111111101111110001111101100001111001"; -- Argumento 522( 3.2029518851052186 Radianes) Función -0.061320736302208245
			 when "1000001011" => Y <= "000000111111101111110001111111100010110011"; -- Argumento 523( 3.2090878082567613 Radianes) Función -0.06744391956366393
			 when "1000001100" => Y <= "000000111111101111110111000111110011011011"; -- Argumento 524( 3.215223731408304 Radianes) Función -0.0735645635996675
			 when "1000001101" => Y <= "000000111111101111110111000111100110011111"; -- Argumento 525( 3.2213596545598464 Radianes) Función -0.07968243797142995
			 when "1000001110" => Y <= "000000111111101111110111111110110111110001"; -- Argumento 526( 3.227495577711389 Radianes) Función -0.08579731234443992
			 when "1000001111" => Y <= "000000111111101111110111001101100001110011"; -- Argumento 527( 3.2336315008629315 Radianes) Función -0.09190895649713252
			 when "1000010000" => Y <= "000000111111101111110111001111111111111110"; -- Argumento 528( 3.2397674240144743 Radianes) Función -0.09801714032956059
			 when "1000010001" => Y <= "000000111111100110000111111001100110110000"; -- Argumento 529( 3.2459033471660166 Radianes) Función -0.10412163387205432
			 when "1000010010" => Y <= "000000111111100110000011000011111101001101"; -- Argumento 530( 3.2520392703175593 Radianes) Función -0.110222207293883
			 when "1000010011" => Y <= "000000111111100110000011000000111111111001"; -- Argumento 531( 3.2581751934691017 Radianes) Función -0.11631863091190446
			 when "1000010100" => Y <= "000000111111100110000100110110011010110011"; -- Argumento 532( 3.2643111166206444 Radianes) Función -0.1224106751992161
			 when "1000010101" => Y <= "000000111111100110000100110111111110110011"; -- Argumento 533( 3.2704470397721868 Radianes) Función -0.12849811079379284
			 when "1000010110" => Y <= "000000111111100110000111100101100111011011"; -- Argumento 534( 3.2765829629237295 Radianes) Función -0.13458070850712606
			 when "1000010111" => Y <= "000000111111100110000011001111111100011111"; -- Argumento 535( 3.2827188860752723 Radianes) Función -0.1406582393328493
			 when "1000011000" => Y <= "000000111111100110000011001100111111110001"; -- Argumento 536( 3.2888548092268146 Radianes) Función -0.14673047445536158
			 when "1000011001" => Y <= "000000111111100110000101101110011011110001"; -- Argumento 537( 3.2949907323783574 Radianes) Función -0.15279718525844346
			 when "1000011010" => Y <= "000000111111100110000101101111111111111111"; -- Argumento 538( 3.3011266555298997 Radianes) Función -0.15885814333386122
			 when "1000011011" => Y <= "000000111111100110000001111101100111110011"; -- Argumento 539( 3.3072625786814425 Radianes) Función -0.16491312048996992
			 when "1000011100" => Y <= "000000111111100110000111000111111101110011"; -- Argumento 540( 3.313398501832985 Radianes) Función -0.17096188876030097
			 when "1000011101" => Y <= "000000111111100110000111000111100011111110"; -- Argumento 541( 3.3195344249845276 Radianes) Función -0.1770042204121487
			 when "1000011110" => Y <= "000000111111100110000111111111110011111110"; -- Argumento 542( 3.32567034813607 Radianes) Función -0.18303988795514067
			 when "1000011111" => Y <= "000000111111100110000111111111100111111110"; -- Argumento 543( 3.3318062712876126 Radianes) Función -0.1890686641498061
			 when "1000100000" => Y <= "000000111111100110000111001110110111111110"; -- Argumento 544( 3.3379421944391554 Radianes) Función -0.19509032201612836
			 when "1000100001" => Y <= "000000111111101001101111111001100000110000"; -- Argumento 545( 3.3440781175906977 Radianes) Función -0.20110463484209176
			 when "1000100010" => Y <= "000000111111101001101111111011100010110000"; -- Argumento 546( 3.3502140407422405 Radianes) Función -0.20711137619221862
			 when "1000100011" => Y <= "000000111111101001101011000011110010110000"; -- Argumento 547( 3.356349963893783 Radianes) Función -0.2131103199160912
			 when "1000100100" => Y <= "000000111111101001101011000011100110110000"; -- Argumento 548( 3.3624858870453256 Radianes) Función -0.21910124015686983
			 when "1000100101" => Y <= "000000111111101001101100110110110111111110"; -- Argumento 549( 3.368621810196868 Radianes) Función -0.2250839113597926
			 when "1000100110" => Y <= "000000111111101001101111100101100001111110"; -- Argumento 550( 3.3747577333484107 Radianes) Función -0.2310581082806711
			 when "1000100111" => Y <= "000000111111101001101111100111100011111110"; -- Argumento 551( 3.380893656499953 Radianes) Función -0.23702360599436695
			 when "1000101000" => Y <= "000000111111101001101011001110011011110011"; -- Argumento 552( 3.3870295796514958 Radianes) Función -0.24298017990326382
			 when "1000101001" => Y <= "000000111111101001101011001111111111110011"; -- Argumento 553( 3.393165502803038 Radianes) Función -0.24892760574571987
			 when "1000101010" => Y <= "000000111111101001101101101101100111111111"; -- Argumento 554( 3.399301425954581 Radianes) Función -0.25486565960451446
			 when "1000101011" => Y <= "000000111111101001101001111111111101110001"; -- Argumento 555( 3.4054373491061236 Radianes) Función -0.2607941179152756
			 when "1000101100" => Y <= "000000111111101001101001111100111111110001"; -- Argumento 556( 3.411573272257666 Radianes) Función -0.26671275747489825
			 when "1000101101" => Y <= "000000111111101001101111000110011010011111"; -- Argumento 557( 3.4177091954092087 Radianes) Función -0.27262135544994903
			 when "1000101110" => Y <= "000000111111101001101111000111111111011011"; -- Argumento 558( 3.423845118560751 Radianes) Función -0.2785196893850529
			 when "1000101111" => Y <= "000000111111101001101111111101100110110011"; -- Argumento 559( 3.429981041712294 Radianes) Función -0.2844075372112719
			 when "1000110000" => Y <= "000000111111101001101111001111111101001101"; -- Argumento 560( 3.436116964863836 Radianes) Función -0.29028467725446216
			 when "1000110001" => Y <= "000000111111101001101111001100111110110000"; -- Argumento 561( 3.442252888015379 Radianes) Función -0.2961508882436238
			 when "1000110010" => Y <= "000000111111101111001111111010011011111110"; -- Argumento 562( 3.448388811166921 Radianes) Función -0.3020059493192278
			 when "1000110011" => Y <= "000000111111101111001111111011100011111111"; -- Argumento 563( 3.454524734318464 Radianes) Función -0.3078496400415348
			 when "1000110100" => Y <= "000000111111101111001011000011110010011111"; -- Argumento 564( 3.4606606574700063 Radianes) Función -0.3136817403988912
			 when "1000110101" => Y <= "000000111111101111001011000011100111011011"; -- Argumento 565( 3.466796580621549 Radianes) Función -0.3195020308160156
			 when "1000110110" => Y <= "000000111111101111001100110110110111111001"; -- Argumento 566( 3.472932503773092 Radianes) Función -0.32531029216226304
			 when "1000110111" => Y <= "000000111111101111001111100101100000110000"; -- Argumento 567( 3.479068426924634 Radianes) Función -0.33110630575987626
			 when "1000111000" => Y <= "000000111111101111001111100100111111111111"; -- Argumento 568( 3.485204350076177 Radianes) Función -0.3368898533922201
			 when "1000111001" => Y <= "000000111111101111001011001110011010011111"; -- Argumento 569( 3.4913402732277192 Radianes) Función -0.3426607173119942
			 when "1000111010" => Y <= "000000111111101111001011001111111110110011"; -- Argumento 570( 3.497476196379262 Radianes) Función -0.34841868024943456
			 when "1000111011" => Y <= "000000111111101111001101101101100110110000"; -- Argumento 571( 3.5036121195308043 Radianes) Función -0.3541635254204902
			 when "1000111100" => Y <= "000000111111101111001101101111100111111111"; -- Argumento 572( 3.509748042682347 Radianes) Función -0.3598950365349881
			 when "1000111101" => Y <= "000000111111101111001001111110110110011111"; -- Argumento 573( 3.5158839658338894 Radianes) Función -0.3656129978047736
			 when "1000111110" => Y <= "000000111111101111001111000101100001111001"; -- Argumento 574( 3.522019888985432 Radianes) Función -0.3713171939518375
			 when "1000111111" => Y <= "000000111111101111001111000111100011111110"; -- Argumento 575( 3.5281558121369745 Radianes) Función -0.3770074102164179
			 when "1001000000" => Y <= "000000111111101111001111111110011010011111"; -- Argumento 576( 3.5342917352885173 Radianes) Función -0.38268343236508967
			 when "1001000001" => Y <= "000000111111101111001111111111111111111001"; -- Argumento 577( 3.54042765844006 Radianes) Función -0.38834504669882636
			 when "1001000010" => Y <= "000000111111101111001111001111110011110011"; -- Argumento 578( 3.5465635815916023 Radianes) Función -0.39399204006104793
			 when "1001000011" => Y <= "000000111111101111001111001111100110011111"; -- Argumento 579( 3.552699504743145 Radianes) Función -0.39962419984564684
			 when "1001000100" => Y <= "000000111111100110011111111010110111001101"; -- Argumento 580( 3.5588354278946874 Radianes) Función -0.4052413140049897
			 when "1001000101" => Y <= "000000111111100110011011000011111101111111"; -- Argumento 581( 3.56497135104623 Radianes) Función -0.4108431710579039
			 when "1001000110" => Y <= "000000111111100110011011000000111110110011"; -- Argumento 582( 3.5711072741977725 Radianes) Función -0.41642956009763693
			 when "1001000111" => Y <= "000000111111100110011100110110011011111110"; -- Argumento 583( 3.5772431973493153 Radianes) Función -0.4220002707997996
			 when "1001001000" => Y <= "000000111111100110011100110111100011011011"; -- Argumento 584( 3.5833791205008576 Radianes) Función -0.4275550934302818
			 when "1001001001" => Y <= "000000111111100110011111100111110011111110"; -- Argumento 585( 3.5895150436524004 Radianes) Función -0.4330938188531519
			 when "1001001010" => Y <= "000000111111100110011111100111111110011111"; -- Argumento 586( 3.5956509668039427 Radianes) Función -0.4386162385385273
			 when "1001001011" => Y <= "000000111111100110011011001101100110110000"; -- Argumento 587( 3.6017868899554855 Radianes) Función -0.4441221445704291
			 when "1001001100" => Y <= "000000111111100110011011001111100110011111"; -- Argumento 588( 3.6079228131070282 Radianes) Función -0.44961132965460665
			 when "1001001101" => Y <= "000000111111100110011101101110110111111110"; -- Argumento 589( 3.6140587362585705 Radianes) Función -0.45508358712634367
			 when "1001001110" => Y <= "000000111111100110011001111111111101011011"; -- Argumento 590( 3.6201946594101133 Radianes) Función -0.46053871095824006
			 when "1001001111" => Y <= "000000111111100110011001111110110111110011"; -- Argumento 591( 3.6263305825616556 Radianes) Función -0.46597649576796596
			 when "1001010000" => Y <= "000000111111100110011111000101100001111001"; -- Argumento 592( 3.6324665057131984 Radianes) Función -0.47139673682599764
			 when "1001010001" => Y <= "000000111111100110011111000100111111110001"; -- Argumento 593( 3.6386024288647407 Radianes) Función -0.4767992300633219
			 when "1001010010" => Y <= "000000111111100110011111111110011010110000"; -- Argumento 594( 3.6447383520162835 Radianes) Función -0.4821837720791227
			 when "1001010011" => Y <= "000000111111100110011111111111100011011011"; -- Argumento 595( 3.650874275167826 Radianes) Función -0.4875501601484357
			 when "1001010100" => Y <= "000000111111100110011111001110011011111111"; -- Argumento 596( 3.6570101983193686 Radianes) Función -0.4928981922297839
			 when "1001010101" => Y <= "000000111111100110011111001111111111001101"; -- Argumento 597( 3.663146121470911 Radianes) Función -0.49822766697278154
			 when "1001010110" => Y <= "000000111111101011011111111011110011011011"; -- Argumento 598( 3.6692820446224537 Radianes) Función -0.5035383837257175
			 when "1001010111" => Y <= "000000111111101011011111111011111111111111"; -- Argumento 599( 3.6754179677739964 Radianes) Función -0.5088301425431071
			 when "1001011000" => Y <= "000000111111101011011011000001100110110000"; -- Argumento 600( 3.6815538909255388 Radianes) Función -0.5141027441932216
			 when "1001011001" => Y <= "000000111111101011011011000011100111111001"; -- Argumento 601( 3.6876898140770815 Radianes) Función -0.5193559901655896
			 when "1001011010" => Y <= "000000111111101011011100110101100111011011"; -- Argumento 602( 3.693825737228624 Radianes) Función -0.5245896826784687
			 when "1001011011" => Y <= "000000111111101011011100110111100111111111"; -- Argumento 603( 3.6999616603801666 Radianes) Función -0.5298036246862946
			 when "1001011100" => Y <= "000000111111101011011111100101100111110011"; -- Argumento 604( 3.706097583531709 Radianes) Función -0.5349976198870969
			 when "1001011101" => Y <= "000000111111101011011011001111111100110000"; -- Argumento 605( 3.7122335066832517 Radianes) Función -0.5401714727298929
			 when "1001011110" => Y <= "000000111111101011011011001110110111111001"; -- Argumento 606( 3.718369429834794 Radianes) Función -0.5453249884220461
			 when "1001011111" => Y <= "000000111111101011011101101111111100110011"; -- Argumento 607( 3.724505352986337 Radianes) Función -0.5504579729366047
			 when "1001100000" => Y <= "000000111111101011011101101110110111011011"; -- Argumento 608( 3.730641276137879 Radianes) Función -0.555570233019602
			 when "1001100001" => Y <= "000000111111101011011001111111111100011111"; -- Argumento 609( 3.736777199289422 Radianes) Función -0.5606615761973359
			 when "1001100010" => Y <= "000000111111101011011001111110110111110001"; -- Argumento 610( 3.7429131224409646 Radianes) Función -0.5657318107836132
			 when "1001100011" => Y <= "000000111111101011011111000111111101110001"; -- Argumento 611( 3.749049045592507 Radianes) Función -0.5707807458869671
			 when "1001100100" => Y <= "000000111111101011011111000110110111111111"; -- Argumento 612( 3.7551849687440497 Radianes) Función -0.5758081914178453
			 when "1001100101" => Y <= "000000111111101011011111111111111101111111"; -- Argumento 613( 3.761320891895592 Radianes) Función -0.5808139580957643
			 when "1001100110" => Y <= "000000111111101011011111111110110111110001"; -- Argumento 614( 3.767456815047135 Radianes) Función -0.5857978574564389
			 when "1001100111" => Y <= "000000111111101011011111001111111101110001"; -- Argumento 615( 3.773592738198677 Radianes) Función -0.590759701858874
			 when "1001101000" => Y <= "000000111111101011011111001110110110011111"; -- Argumento 616( 3.77972866135022 Radianes) Función -0.5956993044924332
			 when "1001101001" => Y <= "000000111111100011111111111011111100011111"; -- Argumento 617( 3.785864584501762 Radianes) Función -0.6006164793838686
			 when "1001101010" => Y <= "000000111111100011111111111010110111011011"; -- Argumento 618( 3.792000507653305 Radianes) Función -0.6055110414043254
			 when "1001101011" => Y <= "000000111111100011111011000011111101111001"; -- Argumento 619( 3.7981364308048478 Radianes) Función -0.6103828062763095
			 when "1001101100" => Y <= "000000111111100011111011000010110111001101"; -- Argumento 620( 3.80427235395639 Radianes) Función -0.6152315905806267
			 when "1001101101" => Y <= "000000111111100011111100110111111101111110"; -- Argumento 621( 3.810408277107933 Radianes) Función -0.6200572117632892
			 when "1001101110" => Y <= "000000111111100011111100110101100111111111"; -- Argumento 622( 3.816544200259475 Radianes) Función -0.6248594881423862
			 when "1001101111" => Y <= "000000111111100011111100110111100110011111"; -- Argumento 623( 3.822680123411018 Radianes) Función -0.629638238914927
			 when "1001110000" => Y <= "000000111111100011111111100101100111111001"; -- Argumento 624( 3.8288160465625602 Radianes) Función -0.6343932841636453
			 when "1001110001" => Y <= "000000111111100011111111100111100110110000"; -- Argumento 625( 3.834951969714103 Radianes) Función -0.6391244448637757
			 when "1001110010" => Y <= "000000111111100011111011001111110011111111"; -- Argumento 626( 3.8410878928656453 Radianes) Función -0.6438315428897913
			 when "1001110011" => Y <= "000000111111100011111011001111111111011011"; -- Argumento 627( 3.847223816017188 Radianes) Función -0.6485144010221124
			 when "1001110100" => Y <= "000000111111100011111101101111110010110000"; -- Argumento 628( 3.8533597391687304 Radianes) Función -0.6531728429537765
			 when "1001110101" => Y <= "000000111111100011111101101111100011111111"; -- Argumento 629( 3.859495662320273 Radianes) Función -0.6578066932970785
			 when "1001110110" => Y <= "000000111111100011111001111110011010110011"; -- Argumento 630( 3.865631585471816 Radianes) Función -0.6624157775901718
			 when "1001110111" => Y <= "000000111111100011111001111100111111110011"; -- Argumento 631( 3.8717675086233583 Radianes) Función -0.6669999223036374
			 when "1001111000" => Y <= "000000111111100011111111000101100001011011"; -- Argumento 632( 3.877903431774901 Radianes) Función -0.6715589548470184
			 when "1001111001" => Y <= "000000111111100011111111000100111111111110"; -- Argumento 633( 3.8840393549264434 Radianes) Función -0.6760927035753158
			 when "1001111010" => Y <= "000000111111100011111111111111111100011111"; -- Argumento 634( 3.890175278077986 Radianes) Función -0.680600997795453
			 when "1001111011" => Y <= "000000111111100011111111111110110111111110"; -- Argumento 635( 3.8963112012295285 Radianes) Función -0.6850836677727002
			 when "1001111100" => Y <= "000000111111100011111111111111100111011011"; -- Argumento 636( 3.902447124381071 Radianes) Función -0.6895405447370669
			 when "1001111101" => Y <= "000000111111100011111111001111110011110011"; -- Argumento 637( 3.9085830475326135 Radianes) Función -0.6939714608896538
			 when "1001111110" => Y <= "000000111111100011111111001111111111111001"; -- Argumento 638( 3.9147189706841563 Radianes) Función -0.6983762494089728
			 when "1001111111" => Y <= "000000111111101110001111111010011011110001"; -- Argumento 639( 3.9208548938356986 Radianes) Función -0.7027547444572251
			 when "1010000000" => Y <= "000000111111101110001111111011100010110000"; -- Argumento 640( 3.9269908169872414 Radianes) Función -0.7071067811865474
			 when "1010000001" => Y <= "000000111111101110001011000001100000110011"; -- Argumento 641( 3.933126740138784 Radianes) Función -0.7114321957452164
			 when "1010000010" => Y <= "000000111111101110001011000010110111110001"; -- Argumento 642( 3.9392626632903265 Radianes) Función -0.7157308252838185
			 when "1010000011" => Y <= "000000111111101110001100110111111101111110"; -- Argumento 643( 3.9453985864418692 Radianes) Función -0.7200025079613817
			 when "1010000100" => Y <= "000000111111101110001100110101100111001101"; -- Argumento 644( 3.9515345095934116 Radianes) Función -0.7242470829514667
			 when "1010000101" => Y <= "000000111111101110001100110111111110110011"; -- Argumento 645( 3.9576704327449543 Radianes) Función -0.7284643904482252
			 when "1010000110" => Y <= "000000111111101110001111100110011010011111"; -- Argumento 646( 3.9638063558964967 Radianes) Función -0.7326542716724126
			 when "1010000111" => Y <= "000000111111101110001111100100111111111111"; -- Argumento 647( 3.9699422790480394 Radianes) Función -0.7368165688773698
			 when "1010001000" => Y <= "000000111111101110001011001111111101110011"; -- Argumento 648( 3.9760782021995817 Radianes) Función -0.7409511253549589
			 when "1010001001" => Y <= "000000111111101110001011001110110111111110"; -- Argumento 649( 3.9822141253511245 Radianes) Función -0.7450577854414658
			 when "1010001010" => Y <= "000000111111101110001011001111100110110000"; -- Argumento 650( 3.988350048502667 Radianes) Función -0.749136394523459
			 when "1010001011" => Y <= "000000111111101110001101101111110010110000"; -- Argumento 651( 3.9944859716542096 Radianes) Función -0.7531867990436123
			 when "1010001100" => Y <= "000000111111101110001101101111100011001101"; -- Argumento 652( 4.000621894805752 Radianes) Función -0.7572088465064842
			 when "1010001101" => Y <= "000000111111101110001001111101100001001101"; -- Argumento 653( 4.006757817957295 Radianes) Función -0.761202385484262
			 when "1010001110" => Y <= "000000111111101110001001111110110110110000"; -- Argumento 654( 4.0128937411088375 Radianes) Función -0.765167265622459
			 when "1010001111" => Y <= "000000111111101110001001111111100110110000"; -- Argumento 655( 4.01902966426038 Radianes) Función -0.7691033376455795
			 when "1010010000" => Y <= "000000111111101110001111000111110011111110"; -- Argumento 656( 4.025165587411922 Radianes) Función -0.7730104533627367
			 when "1010010001" => Y <= "000000111111101110001111000100111111111111"; -- Argumento 657( 4.031301510563465 Radianes) Función -0.7768884656732326
			 when "1010010010" => Y <= "000000111111101110001111111111111101110001"; -- Argumento 658( 4.037437433715008 Radianes) Función -0.7807372285720944
			 when "1010010011" => Y <= "000000111111101110001111111101100111011011"; -- Argumento 659( 4.04357335686655 Radianes) Función -0.784556597155575
			 when "1010010100" => Y <= "000000111111101110001111111111111111111001"; -- Argumento 660( 4.049709280018092 Radianes) Función -0.7883464276266059
			 when "1010010101" => Y <= "000000111111101110001111001110011010110000"; -- Argumento 661( 4.0558452031696355 Radianes) Función -0.7921065773002124
			 when "1010010110" => Y <= "000000111111101110001111001110110111111111"; -- Argumento 662( 4.061981126321178 Radianes) Función -0.7958369046088833
			 when "1010010111" => Y <= "000000111111101110001111001111100111011011"; -- Argumento 663( 4.06811704947272 Radianes) Función -0.7995372691079048
			 when "1010011000" => Y <= "000000111111101111111111111011110011001101"; -- Argumento 664( 4.074252972624263 Radianes) Función -0.803207531480645
			 when "1010011001" => Y <= "000000111111101111111111111000111111111111"; -- Argumento 665( 4.080388895775806 Radianes) Función -0.8068475535437992
			 when "1010011010" => Y <= "000000111111101111111011000011111100110011"; -- Argumento 666( 4.086524818927348 Radianes) Función -0.8104571982525947
			 when "1010011011" => Y <= "000000111111101111111011000001100111111110"; -- Argumento 667( 4.09266074207889 Radianes) Función -0.8140363297059481
			 when "1010011100" => Y <= "000000111111101111111011000011100011011011"; -- Argumento 668( 4.0987966652304335 Radianes) Función -0.8175848131515837
			 when "1010011101" => Y <= "000000111111101111111100110101100000110000"; -- Argumento 669( 4.104932588381976 Radianes) Función -0.8211025149911046
			 when "1010011110" => Y <= "000000111111101111111100110101100111011011"; -- Argumento 670( 4.111068511533518 Radianes) Función -0.8245893027850251
			 when "1010011111" => Y <= "000000111111101111111100110111111111111110"; -- Argumento 671( 4.1172044346850605 Radianes) Función -0.8280450452577554
			 when "1010100000" => Y <= "000000111111101111111111100101100000110011"; -- Argumento 672( 4.123340357836604 Radianes) Función -0.8314696123025452
			 when "1010100001" => Y <= "000000111111101111111111100101100111111111"; -- Argumento 673( 4.129476280988146 Radianes) Función -0.8348628749863799
			 when "1010100010" => Y <= "000000111111101111111111100111111111001101"; -- Argumento 674( 4.135612204139688 Radianes) Función -0.8382247055548377
			 when "1010100011" => Y <= "000000111111101111111011001101100001011011"; -- Argumento 675( 4.1417481272912315 Radianes) Función -0.8415549774368986
			 when "1010100100" => Y <= "000000111111101111111011001101100111111111"; -- Argumento 676( 4.147884050442774 Radianes) Función -0.844853565249707
			 when "1010100101" => Y <= "000000111111101111111011001111111110110000"; -- Argumento 677( 4.154019973594316 Radianes) Función -0.8481203448032971
			 when "1010100110" => Y <= "000000111111101111111101101101100001111001"; -- Argumento 678( 4.1601558967458585 Radianes) Función -0.8513551931052649
			 when "1010100111" => Y <= "000000111111101111111101101101100111011011"; -- Argumento 679( 4.166291819897402 Radianes) Función -0.8545579883654005
			 when "1010101000" => Y <= "000000111111101111111101101111100011110001"; -- Argumento 680( 4.172427743048944 Radianes) Función -0.857728610000272
			 when "1010101001" => Y <= "000000111111101111111001111111111101111111"; -- Argumento 681( 4.178563666200486 Radianes) Función -0.8608669386377671
			 when "1010101010" => Y <= "000000111111101111111001111111110011110011"; -- Argumento 682( 4.184699589352029 Radianes) Función -0.8639728561215865
			 when "1010101011" => Y <= "000000111111101111111001111111100011111110"; -- Argumento 683( 4.190835512503572 Radianes) Función -0.8670462455156926
			 when "1010101100" => Y <= "000000111111101111111111000111111101111110"; -- Argumento 684( 4.196971435655114 Radianes) Función -0.8700869911087113
			 when "1010101101" => Y <= "000000111111101111111111000111110011111110"; -- Argumento 685( 4.2031073588066565 Radianes) Función -0.8730949784182899
			 when "1010101110" => Y <= "000000111111101111111111000100111111111110"; -- Argumento 686( 4.2092432819582 Radianes) Función -0.8760700941954067
			 when "1010101111" => Y <= "000000111111101111111111000111100111111110"; -- Argumento 687( 4.215379205109742 Radianes) Función -0.8790122264286335
			 when "1010110000" => Y <= "000000111111101111111111111101100001110011"; -- Argumento 688( 4.221515128261284 Radianes) Función -0.8819212643483549
			 when "1010110001" => Y <= "000000111111101111111111111101100111110001"; -- Argumento 689( 4.227651051412827 Radianes) Función -0.8847970984309376
			 when "1010110010" => Y <= "000000111111101111111111111111100010011111"; -- Argumento 690( 4.23378697456437 Radianes) Función -0.887639620402854
			 when "1010110011" => Y <= "000000111111101111111111001111111100110011"; -- Argumento 691( 4.239922897715912 Radianes) Función -0.8904487232447579
			 when "1010110100" => Y <= "000000111111101111111111001111110011001101"; -- Argumento 692( 4.246058820867455 Radianes) Función -0.8932243011955152
			 when "1010110101" => Y <= "000000111111101111111111001110110111110011"; -- Argumento 693( 4.252194744018997 Radianes) Función -0.8959662497561849
			 when "1010110110" => Y <= "000000111111101111111111001111111110011111"; -- Argumento 694( 4.25833066717054 Radianes) Función -0.8986744656939538
			 when "1010110111" => Y <= "000000111111101110011111111001100001111001"; -- Argumento 695( 4.264466590322082 Radianes) Función -0.9013488470460219
			 when "1010111000" => Y <= "000000111111101110011111111011110011110011"; -- Argumento 696( 4.270602513473625 Radianes) Función -0.9039892931234431
			 when "1010111001" => Y <= "000000111111101110011111111000111111011011"; -- Argumento 697( 4.276738436625168 Radianes) Función -0.9065957045149154
			 when "1010111010" => Y <= "000000111111101110011111111011100110110000"; -- Argumento 698( 4.28287435977671 Radianes) Función -0.9091679830905224
			 when "1010111011" => Y <= "000000111111101110011011000001100001110001"; -- Argumento 699( 4.289010282928253 Radianes) Función -0.9117060320054298
			 when "1010111100" => Y <= "000000111111101110011011000001100111001101"; -- Argumento 700( 4.295146206079795 Radianes) Función -0.9142097557035305
			 when "1010111101" => Y <= "000000111111101110011011000000111110011111"; -- Argumento 701( 4.301282129231338 Radianes) Función -0.9166790599210427
			 when "1010111110" => Y <= "000000111111101110011011000011100110110000"; -- Argumento 702( 4.3074180523828804 Radianes) Función -0.9191138516900577
			 when "1010111111" => Y <= "000000111111101110011100110101100001011011"; -- Argumento 703( 4.313553975534423 Radianes) Función -0.9215140393420418
			 when "1011000000" => Y <= "000000111111101110011100110111110011111111"; -- Argumento 704( 4.319689898685965 Radianes) Función -0.9238795325112865
			 when "1011000001" => Y <= "000000111111101110011100110100111111001101"; -- Argumento 705( 4.325825821837508 Radianes) Función -0.9262102421383114
			 when "1011000010" => Y <= "000000111111101110011100110111111111011011"; -- Argumento 706( 4.331961744989051 Radianes) Función -0.9285060804732155
			 when "1011000011" => Y <= "000000111111101110011111100111111101110001"; -- Argumento 707( 4.338097668140593 Radianes) Función -0.9307669610789836
			 when "1011000100" => Y <= "000000111111101110011111100110011011110011"; -- Argumento 708( 4.344233591292136 Radianes) Función -0.932992798834739
			 when "1011000101" => Y <= "000000111111101110011111100110110110110000"; -- Argumento 709( 4.3503695144436785 Radianes) Función -0.9351835099389476
			 when "1011000110" => Y <= "000000111111101110011111100111100011111001"; -- Argumento 710( 4.356505437595221 Radianes) Función -0.9373390119125748
			 when "1011000111" => Y <= "000000111111101110011111100111100110110011"; -- Argumento 711( 4.362641360746763 Radianes) Función -0.9394592236021897
			 when "1011001000" => Y <= "000000111111101110011011001101100001011011"; -- Argumento 712( 4.368777283898306 Radianes) Función -0.9415440651830208
			 when "1011001001" => Y <= "000000111111101110011011001111110011011011"; -- Argumento 713( 4.374913207049849 Radianes) Función -0.9435934581619603
			 when "1011001010" => Y <= "000000111111101110011011001110110110011111"; -- Argumento 714( 4.381049130201391 Radianes) Función -0.9456073253805212
			 when "1011001011" => Y <= "000000111111101110011011001111100011011011"; -- Argumento 715( 4.387185053352934 Radianes) Función -0.9475855910177412
			 when "1011001100" => Y <= "000000111111101110011011001111100111011011"; -- Argumento 716( 4.3933209765044765 Radianes) Función -0.9495281805930367
			 when "1011001101" => Y <= "000000111111101110011101101101100000110011"; -- Argumento 717( 4.399456899656019 Radianes) Función -0.9514350209690083
			 when "1011001110" => Y <= "000000111111101110011101101111110011111001"; -- Argumento 718( 4.405592822807561 Radianes) Función -0.9533060403541938
			 when "1011001111" => Y <= "000000111111101110011101101110110110110000"; -- Argumento 719( 4.411728745959104 Radianes) Función -0.9551411683057708
			 when "1011010000" => Y <= "000000111111101110011101101100111111110011"; -- Argumento 720( 4.417864669110647 Radianes) Función -0.9569403357322088
			 when "1011010001" => Y <= "000000111111101110011101101111111111110001"; -- Argumento 721( 4.424000592262189 Radianes) Función -0.9587034748958715
			 when "1011010010" => Y <= "000000111111101110011001111111111100110011"; -- Argumento 722( 4.430136515413731 Radianes) Función -0.9604305194155657
			 when "1011010011" => Y <= "000000111111101110011001111110011010110000"; -- Argumento 723( 4.4362724385652745 Radianes) Función -0.9621214042690416
			 when "1011010100" => Y <= "000000111111101110011001111111110011110001"; -- Argumento 724( 4.442408361716817 Radianes) Función -0.9637760657954398
			 when "1011010101" => Y <= "000000111111101110011001111110110111111001"; -- Argumento 725( 4.448544284868359 Radianes) Función -0.9653944416976893
			 when "1011010110" => Y <= "000000111111101110011001111100111111110011"; -- Argumento 726( 4.454680208019902 Radianes) Función -0.9669764710448522
			 when "1011010111" => Y <= "000000111111101110011001111111111111011011"; -- Argumento 727( 4.460816131171445 Radianes) Función -0.9685220942744174
			 when "1011011000" => Y <= "000000111111101110011111000111111101111110"; -- Argumento 728( 4.466952054322987 Radianes) Función -0.970031253194544
			 when "1011011001" => Y <= "000000111111101110011111000101100001011011"; -- Argumento 729( 4.473087977474529 Radianes) Función -0.9715038909862517
			 when "1011011010" => Y <= "000000111111101110011111000110011011110011"; -- Argumento 730( 4.479223900626073 Radianes) Función -0.9729399522055602
			 when "1011011011" => Y <= "000000111111101110011111000101100111111001"; -- Argumento 731( 4.485359823777615 Radianes) Función -0.9743393827855759
			 when "1011011100" => Y <= "000000111111101110011111000110110111110001"; -- Argumento 732( 4.491495746929157 Radianes) Función -0.9757021300385285
			 when "1011011101" => Y <= "000000111111101110011111000111100011111110"; -- Argumento 733( 4.4976316700806995 Radianes) Función -0.9770281426577543
			 when "1011011110" => Y <= "000000111111101110011111000111111111111001"; -- Argumento 734( 4.503767593232243 Radianes) Función -0.9783173707196277
			 when "1011011111" => Y <= "000000111111101110011111000111100111011011"; -- Argumento 735( 4.509903516383785 Radianes) Función -0.9795697656854405
			 when "1011100000" => Y <= "000000111111101110011111111111111101110001"; -- Argumento 736( 4.516039439535327 Radianes) Función -0.9807852804032303
			 when "1011100001" => Y <= "000000111111101110011111111101100001110011"; -- Argumento 737( 4.522175362686871 Radianes) Función -0.9819638691095554
			 when "1011100010" => Y <= "000000111111101110011111111111110010110000"; -- Argumento 738( 4.528311285838413 Radianes) Función -0.9831054874312163
			 when "1011100011" => Y <= "000000111111101110011111111101100111001101"; -- Argumento 739( 4.534447208989955 Radianes) Función -0.984210092386929
			 when "1011100100" => Y <= "000000111111101110011111111110110111001101"; -- Argumento 740( 4.540583132141498 Radianes) Función -0.9852776423889411
			 when "1011100101" => Y <= "000000111111101110011111111100111111111001"; -- Argumento 741( 4.546719055293041 Radianes) Función -0.9863080972445987
			 when "1011100110" => Y <= "000000111111101110011111111111100011111001"; -- Argumento 742( 4.552854978444583 Radianes) Función -0.9873014181578583
			 when "1011100111" => Y <= "000000111111101110011111111111111111001101"; -- Argumento 743( 4.558990901596125 Radianes) Función -0.9882575677307495
			 when "1011101000" => Y <= "000000111111101110011111111111100110110000"; -- Argumento 744( 4.565126824747668 Radianes) Función -0.9891765099647809
			 when "1011101001" => Y <= "000000111111101110011111001111111101111110"; -- Argumento 745( 4.571262747899211 Radianes) Función -0.9900582102622971
			 when "1011101010" => Y <= "000000111111101110011111001111111101110011"; -- Argumento 746( 4.577398671050753 Radianes) Función -0.99090263542778
			 when "1011101011" => Y <= "000000111111101110011111001101100001110001"; -- Argumento 747( 4.583534594202296 Radianes) Función -0.9917097536690994
			 when "1011101100" => Y <= "000000111111101110011111001110011010110011"; -- Argumento 748( 4.589670517353839 Radianes) Función -0.9924795345987101
			 when "1011101101" => Y <= "000000111111101110011111001111110011001101"; -- Argumento 749( 4.595806440505381 Radianes) Función -0.9932119492347945
			 when "1011101110" => Y <= "000000111111101110011111001111110011110011"; -- Argumento 750( 4.601942363656923 Radianes) Función -0.9939069700023561
			 when "1011101111" => Y <= "000000111111101110011111001101100111011011"; -- Argumento 751( 4.608078286808466 Radianes) Función -0.9945645707342554
			 when "1011110000" => Y <= "000000111111101110011111001110110110110000"; -- Argumento 752( 4.614214209960009 Radianes) Función -0.9951847266721969
			 when "1011110001" => Y <= "000000111111101110011111001110110111110001"; -- Argumento 753( 4.620350133111551 Radianes) Función -0.9957674144676598
			 when "1011110010" => Y <= "000000111111101110011111001100111111111001"; -- Argumento 754( 4.626486056263094 Radianes) Función -0.996312612182778
			 when "1011110011" => Y <= "000000111111101110011111001100111111111111"; -- Argumento 755( 4.632621979414636 Radianes) Función -0.9968202992911657
			 when "1011110100" => Y <= "000000111111101110011111001111100011001101"; -- Argumento 756( 4.638757902566179 Radianes) Función -0.9972904566786902
			 when "1011110101" => Y <= "000000111111101110011111001111100011110001"; -- Argumento 757( 4.6448938257177215 Radianes) Función -0.9977230666441916
			 when "1011110110" => Y <= "000000111111101110011111001111111110110000"; -- Argumento 758( 4.651029748869264 Radianes) Función -0.9981181129001492
			 when "1011110111" => Y <= "000000111111101110011111001111111110110011"; -- Argumento 759( 4.657165672020807 Radianes) Función -0.9984755805732948
			 when "1011111000" => Y <= "000000111111101110011111001111111111110001"; -- Argumento 760( 4.663301595172349 Radianes) Función -0.9987954562051724
			 when "1011111001" => Y <= "000000111111101110011111001111100111111110"; -- Argumento 761( 4.669437518323892 Radianes) Función -0.9990777277526454
			 when "1011111010" => Y <= "000000111111101110011111001111100111111001"; -- Argumento 762( 4.675573441475434 Radianes) Función -0.9993223845883494
			 when "1011111011" => Y <= "000000111111101110011111001111100111011011"; -- Argumento 763( 4.681709364626977 Radianes) Función -0.9995294175010931
			 when "1011111100" => Y <= "000000111111101110011111001111100110011111"; -- Argumento 764( 4.6878452877785195 Radianes) Función -0.9996988186962042
			 when "1011111101" => Y <= "000000111111101110011111001111100111111111"; -- Argumento 765( 4.693981210930062 Radianes) Función -0.9998305817958234
			 when "1011111110" => Y <= "000000111111101110011111001111100111110011"; -- Argumento 766( 4.700117134081604 Radianes) Función -0.9999247018391445
			 when "1011111111" => Y <= "000000111111101110011111001111100111110011"; -- Argumento 767( 4.706253057233147 Radianes) Función -0.9999811752826011
			 when "1100000000" => Y <= "000000100000011111110111111011111101111110"; -- Argumento 768( 4.71238898038469 Radianes) Función -1.0
			 when "1100000001" => Y <= "000000111111101110011111001111100111110011"; -- Argumento 769( 4.718524903536232 Radianes) Función -0.9999811752826011
			 when "1100000010" => Y <= "000000111111101110011111001111100111110011"; -- Argumento 770( 4.724660826687775 Radianes) Función -0.9999247018391445
			 when "1100000011" => Y <= "000000111111101110011111001111100111111111"; -- Argumento 771( 4.7307967498393175 Radianes) Función -0.9998305817958234
			 when "1100000100" => Y <= "000000111111101110011111001111100110011111"; -- Argumento 772( 4.73693267299086 Radianes) Función -0.9996988186962042
			 when "1100000101" => Y <= "000000111111101110011111001111100111011011"; -- Argumento 773( 4.743068596142402 Radianes) Función -0.9995294175010931
			 when "1100000110" => Y <= "000000111111101110011111001111100111111001"; -- Argumento 774( 4.749204519293945 Radianes) Función -0.9993223845883495
			 when "1100000111" => Y <= "000000111111101110011111001111100111111110"; -- Argumento 775( 4.755340442445488 Radianes) Función -0.9990777277526454
			 when "1100001000" => Y <= "000000111111101110011111001111111111110001"; -- Argumento 776( 4.76147636559703 Radianes) Función -0.9987954562051724
			 when "1100001001" => Y <= "000000111111101110011111001111111110110011"; -- Argumento 777( 4.767612288748572 Radianes) Función -0.9984755805732948
			 when "1100001010" => Y <= "000000111111101110011111001111111110110000"; -- Argumento 778( 4.773748211900116 Radianes) Función -0.9981181129001492
			 when "1100001011" => Y <= "000000111111101110011111001111100011110001"; -- Argumento 779( 4.779884135051658 Radianes) Función -0.9977230666441916
			 when "1100001100" => Y <= "000000111111101110011111001111100011001101"; -- Argumento 780( 4.7860200582032 Radianes) Función -0.9972904566786902
			 when "1100001101" => Y <= "000000111111101110011111001100111111111111"; -- Argumento 781( 4.792155981354743 Radianes) Función -0.9968202992911657
			 when "1100001110" => Y <= "000000111111101110011111001100111111111001"; -- Argumento 782( 4.798291904506286 Radianes) Función -0.996312612182778
			 when "1100001111" => Y <= "000000111111101110011111001110110111110001"; -- Argumento 783( 4.804427827657828 Radianes) Función -0.9957674144676598
			 when "1100010000" => Y <= "000000111111101110011111001110110110110000"; -- Argumento 784( 4.81056375080937 Radianes) Función -0.9951847266721969
			 when "1100010001" => Y <= "000000111111101110011111001101100111011011"; -- Argumento 785( 4.816699673960914 Radianes) Función -0.9945645707342554
			 when "1100010010" => Y <= "000000111111101110011111001111110011110011"; -- Argumento 786( 4.822835597112456 Radianes) Función -0.9939069700023561
			 when "1100010011" => Y <= "000000111111101110011111001111110011001101"; -- Argumento 787( 4.828971520263998 Radianes) Función -0.9932119492347946
			 when "1100010100" => Y <= "000000111111101110011111001110011010110011"; -- Argumento 788( 4.8351074434155406 Radianes) Función -0.9924795345987101
			 when "1100010101" => Y <= "000000111111101110011111001101100001110001"; -- Argumento 789( 4.841243366567084 Radianes) Función -0.9917097536690995
			 when "1100010110" => Y <= "000000111111101110011111001111111101110011"; -- Argumento 790( 4.847379289718626 Radianes) Función -0.99090263542778
			 when "1100010111" => Y <= "000000111111101110011111001111111101111110"; -- Argumento 791( 4.853515212870168 Radianes) Función -0.9900582102622971
			 when "1100011000" => Y <= "000000111111101110011111111111100110110000"; -- Argumento 792( 4.859651136021712 Radianes) Función -0.9891765099647809
			 when "1100011001" => Y <= "000000111111101110011111111111111111001101"; -- Argumento 793( 4.865787059173254 Radianes) Función -0.9882575677307495
			 when "1100011010" => Y <= "000000111111101110011111111111100011111001"; -- Argumento 794( 4.871922982324796 Radianes) Función -0.9873014181578584
			 when "1100011011" => Y <= "000000111111101110011111111100111111111001"; -- Argumento 795( 4.878058905476339 Radianes) Función -0.9863080972445988
			 when "1100011100" => Y <= "000000111111101110011111111110110111001101"; -- Argumento 796( 4.884194828627882 Radianes) Función -0.9852776423889412
			 when "1100011101" => Y <= "000000111111101110011111111101100111001101"; -- Argumento 797( 4.890330751779424 Radianes) Función -0.9842100923869291
			 when "1100011110" => Y <= "000000111111101110011111111111110010110000"; -- Argumento 798( 4.896466674930966 Radianes) Función -0.9831054874312164
			 when "1100011111" => Y <= "000000111111101110011111111101100001110011"; -- Argumento 799( 4.902602598082509 Radianes) Función -0.9819638691095554
			 when "1100100000" => Y <= "000000111111101110011111111111111101110001"; -- Argumento 800( 4.908738521234052 Radianes) Función -0.9807852804032304
			 when "1100100001" => Y <= "000000111111101110011111000111100111011011"; -- Argumento 801( 4.914874444385594 Radianes) Función -0.9795697656854406
			 when "1100100010" => Y <= "000000111111101110011111000111111111111001"; -- Argumento 802( 4.921010367537137 Radianes) Función -0.9783173707196278
			 when "1100100011" => Y <= "000000111111101110011111000111100011111110"; -- Argumento 803( 4.92714629068868 Radianes) Función -0.9770281426577543
			 when "1100100100" => Y <= "000000111111101110011111000110110111110001"; -- Argumento 804( 4.933282213840222 Radianes) Función -0.9757021300385286
			 when "1100100101" => Y <= "000000111111101110011111000101100111111001"; -- Argumento 805( 4.9394181369917645 Radianes) Función -0.974339382785576
			 when "1100100110" => Y <= "000000111111101110011111000110011011110011"; -- Argumento 806( 4.945554060143307 Radianes) Función -0.9729399522055603
			 when "1100100111" => Y <= "000000111111101110011111000101100001011011"; -- Argumento 807( 4.95168998329485 Radianes) Función -0.9715038909862518
			 when "1100101000" => Y <= "000000111111101110011111000111111101111110"; -- Argumento 808( 4.957825906446392 Radianes) Función -0.970031253194544
			 when "1100101001" => Y <= "000000111111101110011001111111111111011011"; -- Argumento 809( 4.963961829597935 Radianes) Función -0.9685220942744174
			 when "1100101010" => Y <= "000000111111101110011001111100111111110011"; -- Argumento 810( 4.970097752749477 Radianes) Función -0.9669764710448523
			 when "1100101011" => Y <= "000000111111101110011001111110110111111001"; -- Argumento 811( 4.97623367590102 Radianes) Función -0.9653944416976894
			 when "1100101100" => Y <= "000000111111101110011001111111110011110001"; -- Argumento 812( 4.9823695990525625 Radianes) Función -0.96377606579544
			 when "1100101101" => Y <= "000000111111101110011001111110011010110000"; -- Argumento 813( 4.988505522204105 Radianes) Función -0.9621214042690417
			 when "1100101110" => Y <= "000000111111101110011001111111111100110011"; -- Argumento 814( 4.994641445355648 Radianes) Función -0.9604305194155658
			 when "1100101111" => Y <= "000000111111101110011101101111111111110001"; -- Argumento 815( 5.00077736850719 Radianes) Función -0.9587034748958716
			 when "1100110000" => Y <= "000000111111101110011101101100111111110011"; -- Argumento 816( 5.006913291658733 Radianes) Función -0.9569403357322089
			 when "1100110001" => Y <= "000000111111101110011101101110110110110000"; -- Argumento 817( 5.013049214810275 Radianes) Función -0.9551411683057709
			 when "1100110010" => Y <= "000000111111101110011101101111110011111001"; -- Argumento 818( 5.019185137961818 Radianes) Función -0.9533060403541938
			 when "1100110011" => Y <= "000000111111101110011101101101100000110011"; -- Argumento 819( 5.0253210611133605 Radianes) Función -0.9514350209690084
			 when "1100110100" => Y <= "000000111111101110011011001111100111011011"; -- Argumento 820( 5.031456984264903 Radianes) Función -0.9495281805930368
			 when "1100110101" => Y <= "000000111111101110011011001111100011011011"; -- Argumento 821( 5.037592907416445 Radianes) Función -0.9475855910177413
			 when "1100110110" => Y <= "000000111111101110011011001110110110011111"; -- Argumento 822( 5.043728830567988 Radianes) Función -0.9456073253805213
			 when "1100110111" => Y <= "000000111111101110011011001111110011011011"; -- Argumento 823( 5.049864753719531 Radianes) Función -0.9435934581619604
			 when "1100111000" => Y <= "000000111111101110011011001101100001011011"; -- Argumento 824( 5.056000676871073 Radianes) Función -0.9415440651830209
			 when "1100111001" => Y <= "000000111111101110011111100111100110110011"; -- Argumento 825( 5.062136600022616 Radianes) Función -0.9394592236021898
			 when "1100111010" => Y <= "000000111111101110011111100111100011111001"; -- Argumento 826( 5.0682725231741586 Radianes) Función -0.937339011912575
			 when "1100111011" => Y <= "000000111111101110011111100110110110110000"; -- Argumento 827( 5.074408446325701 Radianes) Función -0.9351835099389477
			 when "1100111100" => Y <= "000000111111101110011111100110011011110011"; -- Argumento 828( 5.080544369477243 Radianes) Función -0.9329927988347391
			 when "1100111101" => Y <= "000000111111101110011111100111111101110001"; -- Argumento 829( 5.086680292628786 Radianes) Función -0.9307669610789837
			 when "1100111110" => Y <= "000000111111101110011100110111111111011011"; -- Argumento 830( 5.092816215780329 Radianes) Función -0.9285060804732156
			 when "1100111111" => Y <= "000000111111101110011100110100111111001101"; -- Argumento 831( 5.098952138931871 Radianes) Función -0.9262102421383115
			 when "1101000000" => Y <= "000000111111101110011100110111110011111111"; -- Argumento 832( 5.105088062083414 Radianes) Función -0.9238795325112866
			 when "1101000001" => Y <= "000000111111101110011100110101100001011011"; -- Argumento 833( 5.111223985234957 Radianes) Función -0.9215140393420419
			 when "1101000010" => Y <= "000000111111101110011011000011100110110000"; -- Argumento 834( 5.117359908386499 Radianes) Función -0.9191138516900579
			 when "1101000011" => Y <= "000000111111101110011011000000111110011111"; -- Argumento 835( 5.123495831538041 Radianes) Función -0.9166790599210428
			 when "1101000100" => Y <= "000000111111101110011011000001100111001101"; -- Argumento 836( 5.129631754689584 Radianes) Función -0.9142097557035306
			 when "1101000101" => Y <= "000000111111101110011011000001100001110001"; -- Argumento 837( 5.135767677841127 Radianes) Función -0.9117060320054299
			 when "1101000110" => Y <= "000000111111101110011111111011100110110000"; -- Argumento 838( 5.141903600992669 Radianes) Función -0.9091679830905225
			 when "1101000111" => Y <= "000000111111101110011111111000111111011011"; -- Argumento 839( 5.148039524144211 Radianes) Función -0.9065957045149156
			 when "1101001000" => Y <= "000000111111101110011111111011110011110011"; -- Argumento 840( 5.154175447295755 Radianes) Función -0.9039892931234433
			 when "1101001001" => Y <= "000000111111101110011111111001100001111001"; -- Argumento 841( 5.160311370447297 Radianes) Función -0.901348847046022
			 when "1101001010" => Y <= "000000111111101111111111001111111110011111"; -- Argumento 842( 5.166447293598839 Radianes) Función -0.898674465693954
			 when "1101001011" => Y <= "000000111111101111111111001110110111110011"; -- Argumento 843( 5.1725832167503825 Radianes) Función -0.895966249756185
			 when "1101001100" => Y <= "000000111111101111111111001111110011001101"; -- Argumento 844( 5.178719139901925 Radianes) Función -0.8932243011955153
			 when "1101001101" => Y <= "000000111111101111111111001111111100110011"; -- Argumento 845( 5.184855063053467 Radianes) Función -0.890448723244758
			 when "1101001110" => Y <= "000000111111101111111111111111100010011111"; -- Argumento 846( 5.190990986205009 Radianes) Función -0.8876396204028542
			 when "1101001111" => Y <= "000000111111101111111111111101100111110001"; -- Argumento 847( 5.197126909356553 Radianes) Función -0.8847970984309377
			 when "1101010000" => Y <= "000000111111101111111111111101100001110011"; -- Argumento 848( 5.203262832508095 Radianes) Función -0.881921264348355
			 when "1101010001" => Y <= "000000111111101111111111000111100111111110"; -- Argumento 849( 5.209398755659637 Radianes) Función -0.8790122264286336
			 when "1101010010" => Y <= "000000111111101111111111000100111111111110"; -- Argumento 850( 5.21553467881118 Radianes) Función -0.8760700941954069
			 when "1101010011" => Y <= "000000111111101111111111000111110011111110"; -- Argumento 851( 5.221670601962723 Radianes) Función -0.8730949784182901
			 when "1101010100" => Y <= "000000111111101111111111000111111101111110"; -- Argumento 852( 5.227806525114265 Radianes) Función -0.8700869911087116
			 when "1101010101" => Y <= "000000111111101111111001111111100011111110"; -- Argumento 853( 5.2339424482658075 Radianes) Función -0.8670462455156929
			 when "1101010110" => Y <= "000000111111101111111001111111110011110011"; -- Argumento 854( 5.240078371417351 Radianes) Función -0.8639728561215866
			 when "1101010111" => Y <= "000000111111101111111001111111111101111111"; -- Argumento 855( 5.246214294568893 Radianes) Función -0.8608669386377673
			 when "1101011000" => Y <= "000000111111101111111101101111100011110001"; -- Argumento 856( 5.252350217720435 Radianes) Función -0.8577286100002722
			 when "1101011001" => Y <= "000000111111101111111101101101100111011011"; -- Argumento 857( 5.258486140871978 Radianes) Función -0.8545579883654008
			 when "1101011010" => Y <= "000000111111101111111101101101100001111001"; -- Argumento 858( 5.264622064023521 Radianes) Función -0.8513551931052651
			 when "1101011011" => Y <= "000000111111101111111011001111111110110000"; -- Argumento 859( 5.270757987175063 Radianes) Función -0.8481203448032973
			 when "1101011100" => Y <= "000000111111101111111011001101100111111111"; -- Argumento 860( 5.2768939103266055 Radianes) Función -0.8448535652497073
			 when "1101011101" => Y <= "000000111111101111111011001101100001011011"; -- Argumento 861( 5.283029833478148 Radianes) Función -0.8415549774368988
			 when "1101011110" => Y <= "000000111111101111111111100111111111001101"; -- Argumento 862( 5.289165756629691 Radianes) Función -0.8382247055548381
			 when "1101011111" => Y <= "000000111111101111111111100101100111111111"; -- Argumento 863( 5.295301679781233 Radianes) Función -0.8348628749863802
			 when "1101100000" => Y <= "000000111111101111111111100101100000110011"; -- Argumento 864( 5.301437602932776 Radianes) Función -0.8314696123025455
			 when "1101100001" => Y <= "000000111111101111111100110111111111111110"; -- Argumento 865( 5.307573526084319 Radianes) Función -0.8280450452577557
			 when "1101100010" => Y <= "000000111111101111111100110101100111011011"; -- Argumento 866( 5.313709449235861 Radianes) Función -0.8245893027850253
			 when "1101100011" => Y <= "000000111111101111111100110101100000110000"; -- Argumento 867( 5.3198453723874035 Radianes) Función -0.8211025149911049
			 when "1101100100" => Y <= "000000111111101111111011000011100011011011"; -- Argumento 868( 5.325981295538946 Radianes) Función -0.817584813151584
			 when "1101100101" => Y <= "000000111111101111111011000001100111111110"; -- Argumento 869( 5.332117218690489 Radianes) Función -0.8140363297059483
			 when "1101100110" => Y <= "000000111111101111111011000011111100110011"; -- Argumento 870( 5.338253141842031 Radianes) Función -0.8104571982525949
			 when "1101100111" => Y <= "000000111111101111111111111000111111111111"; -- Argumento 871( 5.344389064993574 Radianes) Función -0.8068475535437994
			 when "1101101000" => Y <= "000000111111101111111111111011110011001101"; -- Argumento 872( 5.350524988145116 Radianes) Función -0.8032075314806453
			 when "1101101001" => Y <= "000000111111101110001111001111100111011011"; -- Argumento 873( 5.356660911296659 Radianes) Función -0.799537269107905
			 when "1101101010" => Y <= "000000111111101110001111001110110111111111"; -- Argumento 874( 5.3627968344482015 Radianes) Función -0.7958369046088837
			 when "1101101011" => Y <= "000000111111101110001111001110011010110000"; -- Argumento 875( 5.368932757599744 Radianes) Función -0.7921065773002126
			 when "1101101100" => Y <= "000000111111101110001111111111111111111001"; -- Argumento 876( 5.375068680751287 Radianes) Función -0.7883464276266062
			 when "1101101101" => Y <= "000000111111101110001111111101100111011011"; -- Argumento 877( 5.381204603902829 Radianes) Función -0.7845565971555752
			 when "1101101110" => Y <= "000000111111101110001111111111111101110001"; -- Argumento 878( 5.387340527054372 Radianes) Función -0.7807372285720947
			 when "1101101111" => Y <= "000000111111101110001111000100111111111111"; -- Argumento 879( 5.393476450205914 Radianes) Función -0.7768884656732328
			 when "1101110000" => Y <= "000000111111101110001111000111110011111110"; -- Argumento 880( 5.399612373357457 Radianes) Función -0.7730104533627369
			 when "1101110001" => Y <= "000000111111101110001001111111100110110000"; -- Argumento 881( 5.405748296509 Radianes) Función -0.7691033376455797
			 when "1101110010" => Y <= "000000111111101110001001111110110110110000"; -- Argumento 882( 5.411884219660542 Radianes) Función -0.7651672656224592
			 when "1101110011" => Y <= "000000111111101110001001111101100001001101"; -- Argumento 883( 5.418020142812084 Radianes) Función -0.7612023854842622
			 when "1101110100" => Y <= "000000111111101110001101101111100011001101"; -- Argumento 884( 5.424156065963627 Radianes) Función -0.7572088465064846
			 when "1101110101" => Y <= "000000111111101110001101101111110010110000"; -- Argumento 885( 5.43029198911517 Radianes) Función -0.7531867990436126
			 when "1101110110" => Y <= "000000111111101110001011001111100110110000"; -- Argumento 886( 5.436427912266712 Radianes) Función -0.7491363945234597
			 when "1101110111" => Y <= "000000111111101110001011001110110111111110"; -- Argumento 887( 5.442563835418255 Radianes) Función -0.7450577854414658
			 when "1101111000" => Y <= "000000111111101110001011001111111101110011"; -- Argumento 888( 5.448699758569798 Radianes) Función -0.7409511253549592
			 when "1101111001" => Y <= "000000111111101110001111100100111111111111"; -- Argumento 889( 5.45483568172134 Radianes) Función -0.7368165688773701
			 when "1101111010" => Y <= "000000111111101110001111100110011010011111"; -- Argumento 890( 5.460971604872882 Radianes) Función -0.7326542716724133
			 when "1101111011" => Y <= "000000111111101110001100110111111110110011"; -- Argumento 891( 5.4671075280244255 Radianes) Función -0.7284643904482252
			 when "1101111100" => Y <= "000000111111101110001100110101100111001101"; -- Argumento 892( 5.473243451175968 Radianes) Función -0.724247082951467
			 when "1101111101" => Y <= "000000111111101110001100110111111101111110"; -- Argumento 893( 5.47937937432751 Radianes) Función -0.7200025079613819
			 when "1101111110" => Y <= "000000111111101110001011000010110111110001"; -- Argumento 894( 5.485515297479052 Radianes) Función -0.7157308252838191
			 when "1101111111" => Y <= "000000111111101110001011000001100000110011"; -- Argumento 895( 5.491651220630596 Radianes) Función -0.7114321957452164
			 when "1110000000" => Y <= "000000111111101110001111111011100010110000"; -- Argumento 896( 5.497787143782138 Radianes) Función -0.7071067811865477
			 when "1110000001" => Y <= "000000111111101110001111111010011011110001"; -- Argumento 897( 5.50392306693368 Radianes) Función -0.7027547444572256
			 when "1110000010" => Y <= "000000111111100011111111001111111111111001"; -- Argumento 898( 5.5100589900852235 Radianes) Función -0.6983762494089727
			 when "1110000011" => Y <= "000000111111100011111111001111110011110011"; -- Argumento 899( 5.516194913236766 Radianes) Función -0.693971460889654
			 when "1110000100" => Y <= "000000111111100011111111111111100111011011"; -- Argumento 900( 5.522330836388308 Radianes) Función -0.6895405447370672
			 when "1110000101" => Y <= "000000111111100011111111111110110111111110"; -- Argumento 901( 5.5284667595398505 Radianes) Función -0.6850836677727008
			 when "1110000110" => Y <= "000000111111100011111111111111111100011111"; -- Argumento 902( 5.534602682691394 Radianes) Función -0.680600997795453
			 when "1110000111" => Y <= "000000111111100011111111000100111111111110"; -- Argumento 903( 5.540738605842936 Radianes) Función -0.676092703575316
			 when "1110001000" => Y <= "000000111111100011111111000101100001011011"; -- Argumento 904( 5.546874528994478 Radianes) Función -0.6715589548470187
			 when "1110001001" => Y <= "000000111111100011111001111100111111110011"; -- Argumento 905( 5.553010452146021 Radianes) Función -0.6669999223036379
			 when "1110001010" => Y <= "000000111111100011111001111110011010110011"; -- Argumento 906( 5.559146375297564 Radianes) Función -0.6624157775901718
			 when "1110001011" => Y <= "000000111111100011111101101111100011111111"; -- Argumento 907( 5.565282298449106 Radianes) Función -0.6578066932970789
			 when "1110001100" => Y <= "000000111111100011111101101111110010110000"; -- Argumento 908( 5.5714182216006485 Radianes) Función -0.6531728429537771
			 when "1110001101" => Y <= "000000111111100011111011001111111111011011"; -- Argumento 909( 5.577554144752192 Radianes) Función -0.6485144010221123
			 when "1110001110" => Y <= "000000111111100011111011001111110011111111"; -- Argumento 910( 5.583690067903734 Radianes) Función -0.6438315428897915
			 when "1110001111" => Y <= "000000111111100011111111100111100110110000"; -- Argumento 911( 5.589825991055276 Radianes) Función -0.639124444863776
			 when "1110010000" => Y <= "000000111111100011111111100101100111111001"; -- Argumento 912( 5.595961914206819 Radianes) Función -0.6343932841636459
			 when "1110010001" => Y <= "000000111111100011111100110111100110011111"; -- Argumento 913( 5.602097837358362 Radianes) Función -0.629638238914927
			 when "1110010010" => Y <= "000000111111100011111100110101100111111111"; -- Argumento 914( 5.608233760509904 Radianes) Función -0.6248594881423865
			 when "1110010011" => Y <= "000000111111100011111100110111111101111110"; -- Argumento 915( 5.6143696836614465 Radianes) Función -0.6200572117632894
			 when "1110010100" => Y <= "000000111111100011111011000010110111001101"; -- Argumento 916( 5.620505606812989 Radianes) Función -0.6152315905806274
			 when "1110010101" => Y <= "000000111111100011111011000011111101111001"; -- Argumento 917( 5.626641529964532 Radianes) Función -0.6103828062763095
			 when "1110010110" => Y <= "000000111111100011111111111010110111011011"; -- Argumento 918( 5.632777453116074 Radianes) Función -0.6055110414043257
			 when "1110010111" => Y <= "000000111111100011111111111011111100011111"; -- Argumento 919( 5.638913376267617 Radianes) Función -0.6006164793838693
			 when "1110011000" => Y <= "000000111111101011011111001110110110011111"; -- Argumento 920( 5.64504929941916 Radianes) Función -0.5956993044924332
			 when "1110011001" => Y <= "000000111111101011011111001111111101110001"; -- Argumento 921( 5.651185222570702 Radianes) Función -0.5907597018588743
			 when "1110011010" => Y <= "000000111111101011011111111110110111110001"; -- Argumento 922( 5.6573211457222445 Radianes) Función -0.5857978574564391
			 when "1110011011" => Y <= "000000111111101011011111111111111101111111"; -- Argumento 923( 5.663457068873787 Radianes) Función -0.580813958095765
			 when "1110011100" => Y <= "000000111111101011011111000110110111111111"; -- Argumento 924( 5.66959299202533 Radianes) Función -0.5758081914178452
			 when "1110011101" => Y <= "000000111111101011011111000111111101110001"; -- Argumento 925( 5.675728915176872 Radianes) Función -0.5707807458869674
			 when "1110011110" => Y <= "000000111111101011011001111110110111110001"; -- Argumento 926( 5.681864838328415 Radianes) Función -0.5657318107836135
			 when "1110011111" => Y <= "000000111111101011011001111111111100011111"; -- Argumento 927( 5.688000761479957 Radianes) Función -0.5606615761973366
			 when "1110100000" => Y <= "000000111111101011011101101110110111011011"; -- Argumento 928( 5.6941366846315 Radianes) Función -0.5555702330196022
			 when "1110100001" => Y <= "000000111111101011011101101111111100110011"; -- Argumento 929( 5.700272607783043 Radianes) Función -0.550457972936605
			 when "1110100010" => Y <= "000000111111101011011011001110110111111001"; -- Argumento 930( 5.706408530934585 Radianes) Función -0.5453249884220468
			 when "1110100011" => Y <= "000000111111101011011011001111111100110000"; -- Argumento 931( 5.712544454086128 Radianes) Función -0.5401714727298927
			 when "1110100100" => Y <= "000000111111101011011111100101100111110011"; -- Argumento 932( 5.71868037723767 Radianes) Función -0.5349976198870973
			 when "1110100101" => Y <= "000000111111101011011100110111100111111111"; -- Argumento 933( 5.724816300389213 Radianes) Función -0.5298036246862949
			 when "1110100110" => Y <= "000000111111101011011100110101100111011011"; -- Argumento 934( 5.730952223540755 Radianes) Función -0.5245896826784694
			 when "1110100111" => Y <= "000000111111101011011011000011100111111001"; -- Argumento 935( 5.737088146692298 Radianes) Función -0.5193559901655895
			 when "1110101000" => Y <= "000000111111101011011011000001100110110000"; -- Argumento 936( 5.743224069843841 Radianes) Función -0.5141027441932219
			 when "1110101001" => Y <= "000000111111101011011111111011111111111111"; -- Argumento 937( 5.749359992995383 Radianes) Función -0.5088301425431073
			 when "1110101010" => Y <= "000000111111101011011111111011110011011011"; -- Argumento 938( 5.755495916146925 Radianes) Función -0.5035383837257181
			 when "1110101011" => Y <= "000000111111100110011111001111111111001101"; -- Argumento 939( 5.7616318392984684 Radianes) Función -0.49822766697278187
			 when "1110101100" => Y <= "000000111111100110011111001110011011111111"; -- Argumento 940( 5.767767762450011 Radianes) Función -0.49289819222978426
			 when "1110101101" => Y <= "000000111111100110011111111111100011011011"; -- Argumento 941( 5.773903685601553 Radianes) Función -0.4875501601484364
			 when "1110101110" => Y <= "000000111111100110011111111110011010110000"; -- Argumento 942( 5.780039608753096 Radianes) Función -0.4821837720791226
			 when "1110101111" => Y <= "000000111111100110011111000100111111110001"; -- Argumento 943( 5.786175531904639 Radianes) Función -0.4767992300633222
			 when "1110110000" => Y <= "000000111111100110011111000101100001111001"; -- Argumento 944( 5.792311455056181 Radianes) Función -0.4713967368259979
			 when "1110110001" => Y <= "000000111111100110011001111110110111110011"; -- Argumento 945( 5.798447378207723 Radianes) Función -0.4659764957679667
			 when "1110110010" => Y <= "000000111111100110011001111111111101011011"; -- Argumento 946( 5.8045833013592665 Radianes) Función -0.46053871095823995
			 when "1110110011" => Y <= "000000111111100110011101101110110111111110"; -- Argumento 947( 5.810719224510809 Radianes) Función -0.45508358712634395
			 when "1110110100" => Y <= "000000111111100110011011001111100110011111"; -- Argumento 948( 5.816855147662351 Radianes) Función -0.449611329654607
			 when "1110110101" => Y <= "000000111111100110011011001101100110110000"; -- Argumento 949( 5.822991070813893 Radianes) Función -0.4441221445704298
			 when "1110110110" => Y <= "000000111111100110011111100111111110011111"; -- Argumento 950( 5.829126993965437 Radianes) Función -0.43861623853852766
			 when "1110110111" => Y <= "000000111111100110011111100111110011111110"; -- Argumento 951( 5.835262917116979 Radianes) Función -0.4330938188531522
			 when "1110111000" => Y <= "000000111111100110011100110111100011011011"; -- Argumento 952( 5.841398840268521 Radianes) Función -0.42755509343028253
			 when "1110111001" => Y <= "000000111111100110011100110110011011111110"; -- Argumento 953( 5.8475347634200645 Radianes) Función -0.4220002707997995
			 when "1110111010" => Y <= "000000111111100110011011000000111110110011"; -- Argumento 954( 5.853670686571607 Radianes) Función -0.41642956009763726
			 when "1110111011" => Y <= "000000111111100110011011000011111101111111"; -- Argumento 955( 5.859806609723149 Radianes) Función -0.41084317105790424
			 when "1110111100" => Y <= "000000111111100110011111111010110111001101"; -- Argumento 956( 5.8659425328746915 Radianes) Función -0.4052413140049904
			 when "1110111101" => Y <= "000000111111101111001111001111100110011111"; -- Argumento 957( 5.872078456026235 Radianes) Función -0.39962419984564673
			 when "1110111110" => Y <= "000000111111101111001111001111110011110011"; -- Argumento 958( 5.878214379177777 Radianes) Función -0.39399204006104827
			 when "1110111111" => Y <= "000000111111101111001111111111111111111001"; -- Argumento 959( 5.884350302329319 Radianes) Función -0.3883450466988267
			 when "1111000000" => Y <= "000000111111101111001111111110011010011111"; -- Argumento 960( 5.890486225480862 Radianes) Función -0.3826834323650904
			 when "1111000001" => Y <= "000000111111101111001111000111100011111110"; -- Argumento 961( 5.896622148632405 Radianes) Función -0.37700741021641826
			 when "1111000010" => Y <= "000000111111101111001111000101100001111001"; -- Argumento 962( 5.902758071783947 Radianes) Función -0.37131719395183777
			 when "1111000011" => Y <= "000000111111101111001001111110110110011111"; -- Argumento 963( 5.9088939949354895 Radianes) Función -0.36561299780477435
			 when "1111000100" => Y <= "000000111111101111001101101111100111111111"; -- Argumento 964( 5.915029918087033 Radianes) Función -0.359895036534988
			 when "1111000101" => Y <= "000000111111101111001101101101100110110000"; -- Argumento 965( 5.921165841238575 Radianes) Función -0.35416352542049045
			 when "1111000110" => Y <= "000000111111101111001011001111111110110011"; -- Argumento 966( 5.927301764390117 Radianes) Función -0.3484186802494349
			 when "1111000111" => Y <= "000000111111101111001011001110011010011111"; -- Argumento 967( 5.93343768754166 Radianes) Función -0.34266071731199493
			 when "1111001000" => Y <= "000000111111101111001111100100111111111111"; -- Argumento 968( 5.939573610693203 Radianes) Función -0.33688985339222
			 when "1111001001" => Y <= "000000111111101111001111100101100000110000"; -- Argumento 969( 5.945709533844745 Radianes) Función -0.33110630575987654
			 when "1111001010" => Y <= "000000111111101111001100110110110111111001"; -- Argumento 970( 5.9518454569962875 Radianes) Función -0.3253102921622633
			 when "1111001011" => Y <= "000000111111101111001011000011100111011011"; -- Argumento 971( 5.957981380147831 Radianes) Función -0.31950203081601547
			 when "1111001100" => Y <= "000000111111101111001011000011110010011111"; -- Argumento 972( 5.964117303299373 Radianes) Función -0.3136817403988915
			 when "1111001101" => Y <= "000000111111101111001111111011100011111111"; -- Argumento 973( 5.970253226450915 Radianes) Función -0.30784964004153514
			 when "1111001110" => Y <= "000000111111101111001111111010011011111110"; -- Argumento 974( 5.976389149602458 Radianes) Función -0.30200594931922853
			 when "1111001111" => Y <= "000000111111101001101111001100111110110000"; -- Argumento 975( 5.982525072754001 Radianes) Función -0.2961508882436237
			 when "1111010000" => Y <= "000000111111101001101111001111111101001101"; -- Argumento 976( 5.988660995905543 Radianes) Función -0.29028467725446244
			 when "1111010001" => Y <= "000000111111101001101111111101100110110011"; -- Argumento 977( 5.994796919057086 Radianes) Función -0.28440753721127215
			 when "1111010010" => Y <= "000000111111101001101111000111111111011011"; -- Argumento 978( 6.000932842208628 Radianes) Función -0.27851968938505367
			 when "1111010011" => Y <= "000000111111101001101111000110011010011111"; -- Argumento 979( 6.007068765360171 Radianes) Función -0.2726213554499489
			 when "1111010100" => Y <= "000000111111101001101001111100111111110001"; -- Argumento 980( 6.013204688511713 Radianes) Función -0.2667127574748986
			 when "1111010101" => Y <= "000000111111101001101001111111111101110001"; -- Argumento 981( 6.019340611663256 Radianes) Función -0.2607941179152759
			 when "1111010110" => Y <= "000000111111101001101101101101100111111111"; -- Argumento 982( 6.025476534814799 Radianes) Función -0.25486565960451435
			 when "1111010111" => Y <= "000000111111101001101011001111111111110011"; -- Argumento 983( 6.031612457966341 Radianes) Función -0.2489276057457202
			 when "1111011000" => Y <= "000000111111101001101011001110011011110011"; -- Argumento 984( 6.037748381117884 Radianes) Función -0.24298017990326418
			 when "1111011001" => Y <= "000000111111101001101111100111100011111110"; -- Argumento 985( 6.043884304269426 Radianes) Función -0.23702360599436773
			 when "1111011010" => Y <= "000000111111101001101111100101100001111110"; -- Argumento 986( 6.050020227420969 Radianes) Función -0.23105810828067103
			 when "1111011011" => Y <= "000000111111101001101100110110110111111110"; -- Argumento 987( 6.056156150572511 Radianes) Función -0.22508391135979297
			 when "1111011100" => Y <= "000000111111101001101011000011100110110000"; -- Argumento 988( 6.062292073724054 Radianes) Función -0.21910124015687016
			 when "1111011101" => Y <= "000000111111101001101011000011110010110000"; -- Argumento 989( 6.068427996875596 Radianes) Función -0.21311031991609197
			 when "1111011110" => Y <= "000000111111101001101111111011100010110000"; -- Argumento 990( 6.074563920027139 Radianes) Función -0.20711137619221853
			 when "1111011111" => Y <= "000000111111101001101111111001100000110000"; -- Argumento 991( 6.080699843178682 Radianes) Función -0.20110463484209212
			 when "1111100000" => Y <= "000000111111100110000111001110110111111110"; -- Argumento 992( 6.086835766330224 Radianes) Función -0.19509032201612872
			 when "1111100001" => Y <= "000000111111100110000111111111100111111110"; -- Argumento 993( 6.092971689481767 Radianes) Función -0.18906866414980603
			 when "1111100010" => Y <= "000000111111100110000111111111110011111110"; -- Argumento 994( 6.0991076126333095 Radianes) Función -0.18303988795514103
			 when "1111100011" => Y <= "000000111111100110000111000111100011111110"; -- Argumento 995( 6.105243535784852 Radianes) Función -0.17700422041214905
			 when "1111100100" => Y <= "000000111111100110000111000111111101110011"; -- Argumento 996( 6.111379458936394 Radianes) Función -0.17096188876030177
			 when "1111100101" => Y <= "000000111111100110000001111101100111110011"; -- Argumento 997( 6.117515382087937 Radianes) Función -0.16491312048996984
			 when "1111100110" => Y <= "000000111111100110000101101111111111111111"; -- Argumento 998( 6.12365130523948 Radianes) Función -0.15885814333386158
			 when "1111100111" => Y <= "000000111111100110000101101110011011110001"; -- Argumento 999( 6.129787228391022 Radianes) Función -0.15279718525844382
			 when "1111101000" => Y <= "000000111111100110000011001100111111110001"; -- Argumento 1000( 6.135923151542564 Radianes) Función -0.1467304744553624
			 when "1111101001" => Y <= "000000111111100110000011001111111100011111"; -- Argumento 1001( 6.1420590746941075 Radianes) Función -0.1406582393328492
			 when "1111101010" => Y <= "000000111111100110000111100101100111011011"; -- Argumento 1002( 6.14819499784565 Radianes) Función -0.13458070850712642
			 when "1111101011" => Y <= "000000111111100110000100110111111110110011"; -- Argumento 1003( 6.154330920997192 Radianes) Función -0.12849811079379364
			 when "1111101100" => Y <= "000000111111100110000100110110011010110011"; -- Argumento 1004( 6.160466844148735 Radianes) Función -0.12241067519921603
			 when "1111101101" => Y <= "000000111111100110000011000000111111111001"; -- Argumento 1005( 6.166602767300278 Radianes) Función -0.11631863091190484
			 when "1111101110" => Y <= "000000111111100110000011000011111101001101"; -- Argumento 1006( 6.17273869045182 Radianes) Función -0.11022220729388338
			 when "1111101111" => Y <= "000000111111100110000111111001100110110000"; -- Argumento 1007( 6.178874613603362 Radianes) Función -0.10412163387205513
			 when "1111110000" => Y <= "000000111111101111110111001111111111111110"; -- Argumento 1008( 6.1850105367549055 Radianes) Función -0.09801714032956052
			 when "1111110001" => Y <= "000000111111101111110111001101100001110011"; -- Argumento 1009( 6.191146459906448 Radianes) Función -0.09190895649713289
			 when "1111110010" => Y <= "000000111111101111110111111110110111110001"; -- Argumento 1010( 6.19728238305799 Radianes) Función -0.08579731234444028
			 when "1111110011" => Y <= "000000111111101111110111000111100110011111"; -- Argumento 1011( 6.2034183062095325 Radianes) Función -0.07968243797143076
			 when "1111110100" => Y <= "000000111111101111110111000111110011011011"; -- Argumento 1012( 6.209554229361076 Radianes) Función -0.07356456359966743
			 when "1111110101" => Y <= "000000111111101111110001111111100010110011"; -- Argumento 1013( 6.215690152512618 Radianes) Función -0.0674439195636643
			 when "1111110110" => Y <= "000000111111101111110001111101100001111001"; -- Argumento 1014( 6.22182607566416 Radianes) Función -0.06132073630220905
			 when "1111110111" => Y <= "000000111111101111110101101110110110110000"; -- Argumento 1015( 6.227961998815704 Radianes) Función -0.055195244349689775
			 when "1111111000" => Y <= "000000111111101111110011001111100111111110"; -- Argumento 1016( 6.234097921967246 Radianes) Función -0.04906767432741809
			 when "1111111001" => Y <= "000000111111101111110011001110011011110011"; -- Argumento 1017( 6.240233845118788 Radianes) Función -0.04293825693494114
			 when "1111111010" => Y <= "000000111111101111110111100100111111111111"; -- Argumento 1018( 6.2463697682703305 Radianes) Función -0.036807222941359394
			 when "1111111011" => Y <= "000000111111101111110111100111111100011111"; -- Argumento 1019( 6.252505691421874 Radianes) Función -0.030674803176636546
			 when "1111111100" => Y <= "000000111111101111110100110101100111011011"; -- Argumento 1020( 6.258641614573416 Radianes) Función -0.02454122852291245
			 when "1111111101" => Y <= "000000111111101111110011000011111110110011"; -- Argumento 1021( 6.264777537724958 Radianes) Función -0.018406729905805226
			 when "1111111110" => Y <= "000000111111101111110011000010011011001101"; -- Argumento 1022( 6.270913460876501 Radianes) Función -0.012271538285720572
			 when "1111111111" => Y <= "000000111111101111110111111000111110110000"; -- Argumento 1023( 6.277049384028044 Radianes) Función -0.006135884649154477
			 when others => null; 
		 end case; 
	 end process; 
END TABLE; 
